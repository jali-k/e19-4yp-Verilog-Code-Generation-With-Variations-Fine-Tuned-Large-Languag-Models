```
    task Carry4;

        input [1:0] in;
        output [1:0] out;

        begin
            out = in;
            inside = 1;
        end
    endtask