module dff_inst(D, Clock, Resetn, Q);
input D, Clock, Resetn;
output Q;
lpm_ff flipflop(.data(D),.aclr(Resetn),.clock(Clock),.q(Q));
defparam flipflop.lpm_width = 1;
endmodule

module testbench1();
	parameter n = 2;
	reg D;
	reg [n-1:0] a_in = {3'b001, 3'b010};
	reg [n-1:0] b_in = {3'b010, 3'b010};
	reg Clock;
	wire [n-1:0] Q;

	initial begin
	D = 1'b1;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b0;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b1;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b0;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b1;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b0;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b1;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b0;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b1;
	Clock = 0;
	#100;
	Clock = 1;
	#10;
	D = 1'b0;
	Clock = 0;
	#100;