module Prob_7_2_Moore (Detect_Moore