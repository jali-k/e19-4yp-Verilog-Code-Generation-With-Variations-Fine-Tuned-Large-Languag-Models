#### Original Code:
`parameter i`
#### Modifications:
`parameter direction