module tst_wand1(); //testbench
reg [7:0] i1,i2; // Drv1=pull0, Drv2=pull0 -> o = pull0 (wand rule)
wire [7:0] o;
wand1 ww(i1,i2,o);
initial
begin
i1[0] = 0; // Drv1=pull0, Drv2=pull0 -> o = pull0 (wand rule)
i2[0] = 0;
end
initial $monitor($time,"i1=%b,i2=%b,o=%b",i1,i2,o);
initial #8 $stop; // Added stop
endmodule
### Testbench Output:
i1=00000000,i2=00000000,o=00000000
i1=00000000,i2=00000001,o=00000000
i1=00000000,i2=00000010,o=00000000
i1=00000000,i2=00000011,o=00000000
i1=00000000,i2=00000100,o=00000000
i1=00000000,i2=00000101,o=00000000
i1=00000000,i2=00000110,o=00000000
i1=00000000,i2=00000111,o=00000000
i1=00000000,i2=00001000,o=00000000
i1=00000000,i2=00001001,o=00000000
i1=00000000,i2=00001010,o=00000000
i1=00000000,i2=00001011,o=00000000
i1=00000000,i2=00001100,o=00000000
i1=00000000,i2=00001101,o=00000000
i1=00000000,i2=00001110,o=00000000
i1=00000000,i2=00001111,o=00000000
i1=00000000,i2=00010000,o=00000000
i1=00000000,i2=00010001,o=00000000
i1=00000000,i2=00010010,o=00000000
i1=00000000,i2=00010011,o=00000000
i1=00000000,i2=00010100,o=00000000
i1=00000000,i2=00010101,o=00000000
i1=00000000,i2=00010110,o=00000000
i1=00000000,i2=00010111,o=00000000
i1=00000000,i2=00011000,o=00000000
i1=00000000,i2=00011001,o=00000000
i1=00000000,i2=00011010,o=00000000
i1=00000000,i2=00011011,o=00000000
i1=00000000,i2=00011100,o=00000000
i1=00000000,i2=00011101,o=00000000
i1=00000000,i2=00011110,o=00000000
i1=00000000,i2=00011111,o=00000000
i1=00000000,i2=00100000,o=00000000
i1=00000000,i2=00100001,o=00000000
i1=00000000,i2=00100010,o=00000000
i1=00000000,i2=00100011,o=00000000
i1=00000000,i2=00100100,o=00000000
i1=00000000,i2=00100101,o=00000000
i1=00000000,i2=00100110,o=00000000
i1=00000000,i2=00100111,o=00000000
i1=00000000,i2=00101000,o=00000000
i1=00000000,i2=00101001,o=00000000
i1=00000000,i2=00101010,o=00000000
i1=00000000,i2=00101011,o=00000000
i1=00000000,i2=00101100,o=00000000
i1=00000000,i2=00101101,o=00000000
i1=00000000,i2=00101110,o=00000000
i1=00000000,i2=00101111,o=00000000
i1=00000000,i2=00110000,o=00000000
i1=00000000,i2=00110001,o=00000000
i1=00000000,i2=00110010,o=00000000
i1=00000000,i2=00110011,o=00000000
i1=00000000,i2=00110100,o=00000000
i1=00000000,i2=00110101,o=