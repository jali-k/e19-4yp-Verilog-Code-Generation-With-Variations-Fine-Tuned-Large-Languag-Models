// Initializations moved to initial blocks
// Added monitor and stop
// Replaced variable declarations with part-selects, which have been optimized to bit selects.
reg i1,i2;
wire o;