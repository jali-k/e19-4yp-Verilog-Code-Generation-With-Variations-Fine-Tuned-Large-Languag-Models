```
```
### Description of Changes:
```
```

# 05/22/2018 Bugs Fixed
## Test Case 1: Testcase1.v
### Base Verilog Code:
module testbench ();
generate data;
process data;
endmodule
### Variation Instruction:
Add a paramter to the rand module that is used as an input to an internal module inside