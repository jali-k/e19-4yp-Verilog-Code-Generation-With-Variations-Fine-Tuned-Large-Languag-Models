#include <iostream>
using namespace std;

int main()
{
cout << "Hello world!\n";
return 0;
}