module testbench ();
generate struct { rand bit data; } data;
process data;
endmodule
### Expected Output: