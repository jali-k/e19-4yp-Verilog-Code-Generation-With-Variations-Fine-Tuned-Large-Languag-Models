module mux21b (
input wire a,
input wire b,
input wire s,
output reg y // Output must be reg for procedural assignment
);
always @(*)
case (s)
0 : y = a;
1 : y = b;
default: y = 0;
endcase
endmodule
### Simulation Results (a,b,s):
a b s y
00000000000000000000 0 0000000 00000 0000000 0000000
00000000000000000001 1 0000000 00000 0000000 0000000
00000000000000000010 0 0000001 00001 0000000 0000000
00000000000000000011 1 0000001 00001 0000001 0000000
00000000000000000100 0 0000010 00010 0000000 0000000
00000000000000000101 1 0000010 00010 0000011 0000000
00000000000000000110 0 0000011 00011 0000000 0000000
00000000000000000111 1 0000011 00011 0000110 0000000
00000000000000001000 0 0000100 00100 0000000 0000000
00000000000000001001 1 0000100 00100 0000100 0000000
00000000000000001010 0 0000101 00101 0000000 0000000
00000000000000001011 1 0000101 00101 0000101 0000000
00000000000000001100 0 0000110 00110 0000000 0000000
00000000000000001101 1 0000110 00110 0000110 0000000
00000000000000001110 0 0000111 00111 0000000 0000000
00000000000000001111 1 0000111 00111 0000111 0000000
00000000000000010000 0 0001000 01000 0000000 0000000
00000000000000010001 1 0001000 01000 0000100 0000000
00000000000000010010 0 0001001 01001 0000000 0000000
00000000000000010011 1 0001001 01001 0000101 0000000
00000000000000010100 0 0001010 01010 0000000 0000000
00000000000000010101 1 0001010 01010 0000110 0000000
00000000000000010110 0 0001011 01011 0000000 0000000
00000000000000010111 1 0001011 01011 0000111 0000000
00000000000000011000 0 0001100 01100 0000000 0000000
00000000000000011001 1 0001100 01100 0000100 0000000
00000000000000011010 0 0001101 01101 0000000 0000000
00000000000000011011 1 0001101 01101 0000101 0000000
00000000000000011100 0 0001110 01110 0000000 0000000
00000000000000011101 1 0001110 01110 0000110 0000000
00000000000000011110 0 0001111 01111 0000000 0000000
00000000000000011111 1 0001111 01111 0000111 0000000
00000000000000100000 0 0010000 10000 0000000 0000000
00000000000000100001 1 0010000 10000 0000100 0000000
00000000000000100010 0 0010001 10001 0000000 0000000
00000000000000100011 1 0010001 10001 0000101 0000000
00000000000000100100 0 0010010 10010 0000000 00000