module comp
(input wire [N-1:0] x,
input wire [