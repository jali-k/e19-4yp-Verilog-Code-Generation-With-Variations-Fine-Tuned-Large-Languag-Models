class test_gade(
// Inputs
input clk,
input rst_n,

// Outputs
output a,
output a1
);

// Instantiate gade module
gade