module dff_inst(D, Clock, Resetn, Q);
reg D, Resetn, Q;
`