module tst_nor2NOR2NMOS();
  wire a,b,c,d,e,f,g,h,i,j,k,l; // Declare inputs
  wire n_b; // Declare output
  // Instantiate NMOS NOR2
  define gen_block1 nor2NOR2NMOS(.a(a),.b(b),.c(c),.d(d),.e(e