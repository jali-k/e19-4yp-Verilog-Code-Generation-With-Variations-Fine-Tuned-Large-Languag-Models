module reg_8bit; //8-bit register
input [7:0] di; // Data input
input clk; // Clock input
reg [7:0] do; // Data output
always @(posedge clk)
do <= di;
initial
#200 $finish; // Stop simulation endmodule #### 3. Full Adder ##### Base Verilog Code: module add3(//3-bit adder // Input A,B,C. // Output S,C // S = A+B+C, C = 2 bit carry // Input A,B // Output S,C // S = A+B, C = 1 bit carry module add3( input wire a, b, input wire s_in, c_in, output wire s_out, output wire c_out); // Inputs of add3 module // Inputs a,b input wire a,b; // Inputs s_in,c_in input wire s_in,c_in; // Outputs of add3 module // Outputs s_out,c_out output wire s_out,c_out; // Combined inputs, s_in,c_in,a input wire [1:0] s_in,c_in,a; // Combined outputs, s_out,c_out output wire s_out,c_out; // Adder's functionality // Inputs a,b and s_in,c_in assign s_out = a ^ b ^ c_in; assign c_out = (a & b) | (a & c_in) | (b & c_in); endmodule // Instantiation of 3-bit adder module add4( input wire [2:0] a, b, input wire [2:0] s_in, c_in, // Outputs s_out,c_out output wire [2:0] s_out,c_out); // 3 inputs to adder's 3 inputs // 3 outputs from adder's 3 outputs // a,b,s_in,c_in input wire [2:0] a,b,s_in,c_in; // a[2:0],b[2:0],s_in[2:0],c_in[2:0] wire [2:0] s_out,c_out; // s_out[2:0],c_out[2:0] assign s_out[0] = a[0]^b[0]; assign s_out[1] = a[0]^b[1]^c_in[0]; assign s_out[2] = a[1]^b[1]^c_in[1]; assign c_out[0] = s_in[0]^a[1]^b[0]; assign c_out[1] = s_in[1]^a[1]^b[1]; assign c_out[2] = c_in[1]; endmodule // Instantiation of 4-bit adder module add3( input wire a, b, input wire s_in, c_in, output wire s_out, output wire c_out); add4 add1(.a(a),.b(b),.s_in(s_in),.c_in(c_in),.s_out(s_out),.c_out(c_out)); endmodule // Instantiation of 3-bit adder module add3( input wire a, b, input wire s_in, c_in, output wire s_out, output wire c_out); add4 add1(.a(a),.b(b),.s_in(s_in),.c_in(c_in),.s_out(s_out),.c_out(c_out)); endmodule ##### Variation Instruction: Add `inside` operator to check `s_cnt` inside a constant array and wrap combinational block in escaped generate block. ##### Modified Code: module add3( //3-bit adder // Input A,B,C // Output S,C // S = A+B+C, C = 2 bit carry // Input A,B input wire a,b; // Inputs s_in,c_in input wire s_in,c_in; // Outputs of add3 module // Outputs s_out,c_out output wire s_out,c_out; // Combined inputs, s_in,c_in,a input wire [1:0] s_in,c_in,a; // Combined outputs, s_out,c_out output wire s_out,c_out; // Adder's functionality // Inputs a,b and s_in,c_in assign s_out = a ^ b ^ c_in; assign c_out = (a & b) | (a & c_in) | (b & c_in); endmodule // Instantiation of 3-bit adder module add4( input wire [2:0] a, b, input wire [2:0] s_in, c_in, // Outputs s_out,c_out output wire [2:0] s_out,c_out); // 3 inputs to adder's 3 inputs // 3 outputs from adder's 3 outputs // a,b,s_in,c_in input wire [2:0] a,b,s_in,c_in; // a[2:0],b[2:0],s_in[2:0],c_in[2:0] wire [2:0] s_out,c_out; // s_out[2:0],c_out[2:0] assign s_out[0] = a[0]^b[0]; assign s_out[1] = a[0]^b[1]^c_in[0]; assign s_out[2] = a[1]^b[1]^c_in[1]; assign c_out[0] = s_in[0]^a[1]^b[0]; assign c_out[1] = s_in[1]^a[1]^b[1]; assign c_out[2] = c_in[1]; endmodule // Instantiation of 4-bit adder module add3( input wire a, b, input wire s_in, c_in, output wire s_out, output wire c_out); add4 add1(.a(a),.b(b),.s_in(s_in),.c_in(c_in),.s_out(s_out),.c_out(c_out)); endmodule // Instantiation of 3-bit adder module add3( input wire a, b, input wire s_in, c_in, output wire s_out, output wire c_out); add4 add1(.a(a),.b(b),.s_in(s_in),.c_in(c_in),.s_out(s_out),.c_out(c_out)); endmodule ##### Variation Instruction: Add `inside` operator to check `s_cnt` inside a constant array and wrap combinational block in escaped generate block. ##### Modified Code: module add3( //3-bit adder // Input A,B,C // Output S,C // S = A+B+C, C = 2 bit carry // Input A,B input wire a,b; // Inputs s_in,c_in input wire s_in,c_in; // Outputs of add3 module // Outputs s_out,c_out output wire s_out,c_out; // Combined inputs, s