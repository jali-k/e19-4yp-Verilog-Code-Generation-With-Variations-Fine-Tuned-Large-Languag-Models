module mux41b (
input wire [3:0] c,
input wire [1:0] s,
output wire z
);
wire c1,c2,c3,c4; // Testing array elements
assign {c1,c2} = c[2:0]; // Testing array elements
assign {c3,c4} = c[3:0]; // Testing array elements
case (s)
3'h0: z = ~s[1] & ~s[0] & c[0];
3'h1: z = ~s[1] & s[0] & c[1];
3'h2: z = s[1] & ~s[0] & c2;
3'h3: z = s[1] & s[0] & c3;
default: z = s[1] & s[0] & c4;
endcase
endmodule
### Output:
1) Mux41b:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
2) Mux41b_2:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
3) Mux41b_3:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
4) Mux41b_2_2:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
5) Mux41b_3_2:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
6) Mux41b_3_3:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
7) Mux41b_3_4:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
8) Mux41b_3_5:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
9) Mux41b_3_6:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
10) Mux41b_3_7:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
11) Mux41b_3_8:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3
12) Mux41b_3_9:
1 0 0 1 1 0 0 1 1 0 0 1 1 0 0 1
0 1 2 3 3 3 3 3 3 3 3 3 3 3 3 3