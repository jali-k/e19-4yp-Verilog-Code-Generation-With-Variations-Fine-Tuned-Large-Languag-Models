module Problem2(input [3:0] a, b);
endmodule
module Problem