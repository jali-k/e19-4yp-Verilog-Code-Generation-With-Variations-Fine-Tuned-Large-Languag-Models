/**
 * File Name: ttst_ttrimux2_1.v
 * Designer : Amir Malekpour
 * Date	: Sat May 16 16:04:39 2020
 * Description:
 * 	This is a testbench for tristate 2-to-1 mux.
 * 	Verilog language variant : SystemVerilog
 */
module ttst_ttrimux2_1(); // Assuming this tests a tristate 2-to-1 mux called ttrimux2_1
reg e;
reg [1:0]i; // Should be reg i0, i1; or reg [0:0] i0, i1; or just input wires if MUX takes separate inputs
reg s;
wire out; // Added wire declaration
// ttrimux2_1 mm(out,e,i,s); // Instantiation requires correct MUX definition
initial
begin
e =0; i = 2'b00; s = 1'b0; // Added initial's'