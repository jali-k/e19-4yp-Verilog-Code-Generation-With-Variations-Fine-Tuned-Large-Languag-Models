module AND_test;
reg [3:0] a;
wire [0:0]b;
always @(a)
begin
if (a[3: