Verilog code for