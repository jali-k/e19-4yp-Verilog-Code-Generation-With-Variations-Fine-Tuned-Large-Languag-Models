enum {RESET,SET} Resetn;