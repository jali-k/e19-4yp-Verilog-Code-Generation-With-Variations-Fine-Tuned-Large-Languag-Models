struct packed {
  signed [1:0] a;
  signed [1:0] b;
};
module fa_1(d,s,ci);
  packed {
    a,b} p_in;
  packed {
    d,s} p_out;
  xor #(p_in.a,p_in.b,d);
  and #(p_in.a,p_in.b,ci,s);
endmodule
### Testbench Code:
module tb_fa_1;
  reg a,b;
  wire [1:0] d;
  wire [1:0] s;
  wire [1:0] ci;
  fa_1 inst
  (.d(d),.s(s),.ci(ci),.a(a),.b(b));
  initial $monitor("d=%0h, s=%0h, ci=%0h", d, s, ci);
  initial begin
    repeat(5) begin
      a = 0;
      b = 0;
      #1 a = 1; #1 b = 1; #1 ci = 1;
      #1 a = 0; #1 b = 1; #1 ci = 0;
      #1 a = 1; #1 b = 0; #1 ci = 1;
      #1 a = 0; #1 b = 0; #1 ci = 0;
    end
    $finish;
  end
endmodule
### Wavedrom Source:
#Title: Full Adder
#Author: 
#Generated by: 
#Source: https://www.wavedrom.com/
{signal: [
    {name: "a", wave: "0"},
    {name: "b", wave: "0.1"},
    {name: "ci", wave: "0"},
    {name: "d", wave: "0"},
    {name: "s", wave: "0"}
  ],
  head: {
    text: "Full Adder",
    left: "a",
    right: "b"
  },
  body: [
    {
      head: {
        text: "d",
        left: "a",
        right: "b"
      },
      body: [
        {
          text: "xor (a, b, d)",
          top: "d",
          bottom: "a",
          right: "b"
        },
        {
          text: "and (a, b, ci, s)",
          right: "ci",
          top: "d",
          bottom: "a"
        }
      ]
    }
  ]
}
### Results:
#### Wavedrom:
![wavedrom_fa_1.svg](https://github.com/hawkin8