module example16(clk, rst, q);
input clk, rst;
output