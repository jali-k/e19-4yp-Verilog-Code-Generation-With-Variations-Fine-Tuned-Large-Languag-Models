module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
reg[3:0] a1,b1;
logic[3