```verilog
module reg4_condition(D, Clock, Resetn, Q);
input [3:0] D;
input Clock, Reset