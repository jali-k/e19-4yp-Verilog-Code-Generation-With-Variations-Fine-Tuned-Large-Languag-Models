We will use the same array slice defined in the package:
```verilog
import mixed_sim_