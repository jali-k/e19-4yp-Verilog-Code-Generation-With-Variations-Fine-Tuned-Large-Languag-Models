module example3(Data