module SchedDelayA;
class Sched;
endclass
reg a, b;
initial
begin
end
always b = (Sched)b;
always a = (Sched)b;
endmodule