module dffen(output do,input di,input en);// Instantiate the D latch
reg [3:0] s_cnt = 0;
generate// Generate block
// Add `inside` operator to check `s_cnt` inside a constant array and wrap combinational block in escaped generate block.
for (s_cnt inside {0,1,2,3}) begin
if (en==1) do=di; // if enable is high, then data input is the data output
end
endgenerate// end generate block
endmodule
### Test Output:

en=0, di=0, do=0
en=1, di=0, do=0
en=1, di=1, do=1
en=1, di=0, do=1
en=1, di=0, do=0
en=1, di=0, do=1
en=1, di=1, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=1, di=1, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=1, di=1, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=1, di=1, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=1, di=1, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=1, di=1, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=1, di=1, do=1
en=1, di=0, do=1
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=1, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=0, di=0, do=0
en=