module Prob_13 (Nand_2, di