module VMP_FIFO
(
output [7:0] Data,
output [3:0] Ena,
input  [2:0] Clk,
input  [7:0] WData,
input  [3:0] WEna
);
endmodule

## 3.566.1