module example3(Data, Clock, Reset, RegSum, Sum, ld);
input Clock, Reset;
input [3:0] Data;
output