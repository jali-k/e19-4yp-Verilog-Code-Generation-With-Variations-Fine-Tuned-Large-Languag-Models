module aoi2(g,a,b,c,d);
output g;
input a,b,c,d