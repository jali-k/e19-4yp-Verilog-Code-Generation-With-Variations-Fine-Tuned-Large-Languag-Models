module mux4_4(in[3:0], sel, out);
input [3:0]