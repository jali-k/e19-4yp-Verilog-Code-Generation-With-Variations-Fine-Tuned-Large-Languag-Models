{% set params={ 'clk','N','En' } %}
{% include 'inside_range.v' %}
### Output:
{% set params={ 'clk','N','En' } %}
{% include 'inside_range.v.log' %}