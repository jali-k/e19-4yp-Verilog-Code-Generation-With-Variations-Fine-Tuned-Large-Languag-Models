#### Variation:
```
interface if_a #(parameter p=4)(); // modified to add parameter
logic