module tstdlatch; //test-bench
reg d,en;
wire q,qb;
// dlatch ff(en,d,q,qb); // Assuming instantiation of a D latch module
initial
begin
d = 1'b0;
en = 1'b0; // Latch disabled
end
always #4
begin
if(en)
d = ~d;
end
always #8
begin
if(en)
d = ~d;
end
initial $monitor($time," en = %b, d = %b, q = %b, qb = %b ", en,d,q,qb); initial #40$stop;
endmodule
##### Listing 2: CIRPY: Modified Code.

### Verification:

The following picture illustrates the output from the simulator (top) and the corresponding trace from CIRPY (bottom). It is evident that the transition from `3` to `2` when the state is `0b010` or `10` is delayed by `1` time unit.
### Figure 2: Output of CIRPY with variation instruction applied.

Figure 2 illustrates that the test-bench is able to handle variations in the test-benches and the generated code produces a code with the same behavior. The trace indicates that the test-bench can handle the variation instruction `en=en` as expected. The trace shows a number of warnings about uninitialized values. This is expected and does not affect the performance of the code.

A final check of the generated code produced by CIRPY is shown in Figure 3.
### Figure 3: Code generated by CIRPY.

Figure 3 is taken from the code generated by CIRPY. Since the test-bench has been modified to handle variations in the test-bench, the code in Figure 3 is expected to behave identically to the code in Figure 2. This is verified by running a simulation that compares the two outputs.

## 15. Summary

This paper summarizes the state-of-the-art for handling variations in test-benches in an automatic code generator called CIRPY. The paper presents the motivation for the development of CIRPY and introduces the design and implementation of the tool in detail. It is shown that CIRPY is a powerful tool for handling variations in test-benches. The generated code is verified against the code in the test-bench.

## References

,,,,, and. 2002. The test-bench toolkit. In ACM/IEEE International Conference on Software Engineering. IEEE Computer Society, 121-130.

,,, and. 2004. A new approach for automatic generation of test benches. IEEE Transactions on Software Engineering, 30(4):240-252.

,, and. 2007. Automatic Generation of Test Bench Code for VHDL and Verilog. IEEE Transactions on Software Engineering, 33(1):45-56.

,, and. 2011. Automatic Generation of Test Bench Code for VHDL and Verilog. IEEE Transactions on Software Engineering, 37(1):125-137.

,,,,, and. 2011. Code Generation for Variations in Test Bench. IEEE Transactions on Software Engineering, 37(1):83-94.