module muxdff(D0, D1, Sel, Clock, Q);
input D0, D1, Sel, Clock;
output Q;
reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D0;
    else
        Q <= D1;
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module muxdff(D[0], D[1], Sel, Clock, Q);
input [1:0] D;
input Sel, Clock;
output reg Q;
always @(posedge Clock)
    if (!Sel)
        Q <= D[0];
    else
        Q <= D[1];
endmodule

module m