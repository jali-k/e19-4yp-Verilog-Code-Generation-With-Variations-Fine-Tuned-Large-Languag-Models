module Test (inout a, inout b, inout c);
(a -> b) =