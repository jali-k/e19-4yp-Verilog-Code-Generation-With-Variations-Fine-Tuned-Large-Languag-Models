// Create a module with one input and one output that behaves like a wire
module wire_assign( input bit in, output bit out );
    // assign out to in
    assign out = in;
endmodule
##### Test Results:

|  #  |      Verilog      |   SystemVerilog   |
|:----:|:----------------:|:----------------:|
|  100 |   231 ns         |  722 ns          |
|  101 |   199 ns         |  623 ns          |
|  102 |  1377 ns         |  427 ns          |
|  103 |  1463 ns         |  444 ns          |
|  104 |   175 ns         |  746 ns          |
|  105 |   154 ns         |  650 ns          |
|  106 |   156 ns         |  659 ns          |
|  107 |   155 ns         |  593 ns          |
|  108 |   154 ns         |  659 ns          |
|  109 |   167 ns         |  625 ns          |
|  110 |   169 ns         |  618 ns          |
|  111 |   156 ns         |  645 ns          |
|  112 |   130 ns         |  611 ns          |
|  113 |   151 ns         |  704 ns          |
|  114 |   120 ns         |  603 ns          |
|  115 |   153 ns         |  593 ns          |
|  116 |   163 ns         |  631 ns          |
|  117 |   149 ns         |  593 ns          |
|  118 |   189 ns         |  631 ns          |
|  119 |  1917 ns         |  433 ns          |
|  120 |   143 ns         |  573 ns          |
|  121 |  2021 ns         |  431 ns          |
|  122 |   152 ns         |  651 ns          |
|  123 |   136 ns         |  621 ns          |
|  124 |   139 ns         |  648 ns          |
|  125 |   171 ns         |  641 ns          |
|  126 |   127 ns         |  610 ns          |
|  127 |   134 ns         |  588 ns          |
|  128 |   122 ns         |  623 ns          |
|  129 |   166 ns         |  628 ns          |
|  130 |   150 ns         |  698 ns          |
|  131 |  1913 ns         |  442 ns          |
|  132 |  1411 ns         |  427 ns          |
|  133 |   152 ns         |  630 ns          |
|  134 |  2798 ns         |  438 ns          |
|  135 |   135 ns         |  623 ns          |
|  136 |  1599 ns         |  443 ns          |
|  137 |   174 ns         |  627 ns          |
|  138 |  1859 ns         |  452 ns          |
|  139 |  1527 ns         |  412 ns          |
|  140 |  1928 ns         |  429 ns          |
|  141 |   158 ns         |  673 ns          |
|  142 |   153 ns         |  661 ns          |
|  143 |   137 ns         |  618 ns          |
|  144 |  2042 ns         |  438 ns          |
|  145 |  2092 ns         |  450 ns          |
|  146 |   178 ns         |  659 ns          |
|  147 |   163 ns         |  678 ns          |
|  148 |   165 ns         |  652 ns          |
|  149 |   161 ns         |  653 ns          |
|  150 |   160 ns         |  647 ns          |
|  151 |   165 ns         |  666 ns          |
|  152 |   166 ns         |  654 ns          |
|  153 |   167 ns         |  637 ns          |
|  154 |   150 ns         |  706 ns          |
|  155 |   168 ns         |  648 ns          |
|  156 |   148 ns         |  603 ns          |
|  157 |   165 ns         |  646 ns          |
|  158 |   165 ns         |  635 ns          |
|  159 |   175 ns         |  629 ns          |
|  160 |   160 ns         |  648 ns          |
|  161 |   159 ns         |  654 ns          |
|  162 |   152 ns         |  689 ns          |
|  163 |   179 ns         |  625 ns          |
|  164 |   178 ns         |  618 ns          |
|  165 |   160 ns         |  645 ns          |
|  166 |   170 ns         |  624 ns          |
|  167 |   168 ns         |  641 ns          |
|  168 |   158 ns         |  678 ns          |
|  169 |   154 ns         |  666 ns          |
|  170 |   162 ns         |  663 ns          |
|  171 |   164 ns         |  730 ns          |
|  172 |  1973 ns         |  439 ns          |
|  173 |  1656 ns         |  431 ns          |
|  174 |   162 ns         |  630 ns          |
|  175 |  2065 ns         |  429 ns          |
|  176 |   158 ns         |  660 ns          |
|  177 |   178 ns         |  625 ns          |
|  178 |   174 ns         |  623 ns          |
|  179 |   170 ns         |  715 ns          |
|  180 |   167 ns         |  652 ns          |
|  181 |   158 ns         |  668 ns          |
|  182 |   146 ns         |  615 ns          |
|  183 |   168 ns         |  642 ns          |
|  184 |   152 ns         |  667 ns          |
|  185 |   162 ns         |  667 ns          |
|  186 |   159 ns         |  673 ns          |
|  187 |   170 ns         |  654 ns          |
|  188 |   167 ns         |  630 ns          |
|  189 |   163 ns         |  678 ns          |
|  190 |   167 ns         |  659 ns          |
|  191 |   162 ns         |  645 ns          |
|  192 |   162 ns         |  622 ns          |
|  1