module tb_TOP7;
  reg CLK, RST