`inside` on `state_Moore`