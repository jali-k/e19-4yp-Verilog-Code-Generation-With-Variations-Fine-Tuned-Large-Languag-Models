module testbench ();
generate
struct { rand bit a; } my_data;
endgenerate
process data;
endmodule