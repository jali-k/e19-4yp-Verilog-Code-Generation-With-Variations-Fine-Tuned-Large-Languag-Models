sudo apt-get install socfpga-sw