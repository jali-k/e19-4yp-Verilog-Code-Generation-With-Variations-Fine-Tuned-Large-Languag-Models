module Universal_Shift_Reg (Data_Out, MSB_Out, LSB_Out, Data_In,
MSB_In, LSB_In, s1, s0, clk, rst);
output [3: 0] Data_Out;
output MSB_Out, LSB_Out;
input [3: 0] Data_In;
input MSB_In, LSB_In;
reg [3: 0] Data_Out; // 10-12-2004
input s1, s0, clk, rst;
assign MSB_Out = Data_Out[3];
assign LSB_Out = Data_Out[0];
always @ (posedge clk) begin
if (rst) Data_Out <= 0;
else case (s1, s0)
(0, 0): Data_Out <= Data_Out; // Idle
(.T..T): Data_Out <= {MSB_In, Data_Out[3:1]}; // Shift right
(0,.T): Data_Out <= {Data_Out[2:0], LSB_In}; // Shift Left
(.T, 0): Data_Out <= Data_In; // Parallel Load
(.T,.T): Data_Out <= Data_Out; // reset-on-the-fly
endcase
end
endmodule
/*
Test Plan
Verify initial reset
Verify idle
Verify shift right
Verify shift left
Verify parallel load
Verify reset-on-the-fly
*/
module t_Universal_Shift_Reg();
wire [3: 0] Data_Out;
reg [3: 0] Data_In;
wire MSB_Out, LSB_Out;
reg MSB_In, LSB_In;
reg s1, s0, rst;
defparam M2.half_cycle = 5;

Universal_Shift_Reg M1 (Data_Out, MSB_Out, LSB_Out, Data_In, MSB_In, LSB_In, s1,
s0, clk, rst);
Clock_Gen M2(clk);

initial #1000 $finish;
initial fork
begin #5 rst = 1; #20 rst = 0;end
begin #120 rst = 1; #20 rst = 0;end
begin #260 rst = 1; #20 rst = 0;end
begin #380 rst = 1; #20 rst = 0;end
join
initial fork
join
begin // Verify left shift
join
begin // Verify load
join
begin // reset
join
module Clock_Gen(clk, half_cycle);
input clk;
defparam half_cycle = 5;
output reg clk;
reg half_cycle;
always #half_cycle clk = ~clk;
endmodule
endmodule

## Tips for writing testbenches with VeriLog

### How to write a testbench

The testbench will mostly contain the following tasks:

• A module that needs to be tested
• An instance of the module being tested
• A Clock generator using the defparam system task
• The $finish task
• A reset state
• The testbenches should start with an initial fork that creates all the necessary objects.
• The fork task should contain all the objects that are not needed in the test.
• The initial task should contain any other necessary things, like a reset signal and a $finish task.
• The fork task should contain all the individual tasks that the testbench needs. The tasks can be written out, but it is often better to wrap them in an initial task so that they can be started at the same time.

The individual testbenches should follow a similar structure. There are a few common components.

#### Common Components

The following components will be used across most of the testbenches. In this section, the components will be explained and also the testbenches will be explained. It is recommended to have one testbench per component so that the components can be easily reused in future testbenches.

• Clock Generator:
The clock generator is used to test a clocked module. This can be used to test the reset as well. The testbench will also require a reset signal which will be used to determine the initial state of the module.

The clock generator is used to generate a clock signal. It can be used to test a clocked module and also to test a reset signal. The clock signal is generated using the following code:

module Clock_Gen(clk, half_cycle);
input clk;
defparam half_cycle = 5;
output reg clk;
reg half_cycle;
always #half_cycle clk = ~clk;
endmodule

The clock generator has a clock signal and half_cycle parameter. The clock signal is the clock that is generated by the clock generator. This can be used to test a clocked module. The default value for half_cycle is 5. As the clock signal is generated using the code, the half_cycle parameter is used to decide the period of the clock signal. For example, if the half_cycle is 5 then the clock signal is generated every 5ns. The output clk is generated using the code. The output clk is a register in the code and it is assigned a value using the following code:

reg half_cycle;
always #half_cycle clk = ~clk;

clk is the signal that is generated using the system task. It is assigned the opposite value of the clk signal. This ensures that after every clock edge, the clk signal will have the opposite value. The half_cycle parameter is used to ensure that the clock signal is generated at the proper speed.

• Reset:

The reset task is an optional task that is used to set the reset signal. The reset signal is used to determine the initial state of the module being tested. This is particularly useful for clocked modules. The task is written as follows:

initial fork
begin // Reset the module
initial rst = 1; // Assert the reset signal
join
initial rst = 0; // De-assert the reset signal
join;

This task will assert the reset signal, de-assert it after 5 cycles and then assert it after 25ns.

• Testbench:

The testbench is the actual executable code written in Verilog. The testbenches should start with an initial fork that creates all the necessary objects. The fork should contain all the objects that are not needed in the test. The initial task should contain any other necessary things, like a reset signal and a $finish task. The fork task should contain all the individual tasks that the testbench needs. The tasks can be written out, but it is often better to wrap them in an initial task so that they can be started at the same time. The individual tasks are as follows: 1. The input variables are connected to the corresponding output variables that are being tested: module testbench(); input [3: 0] Data_Out; output [3: 0] Data_In; initial begin fork join initial Data_In = 0; join end fork join endmodule  This testbench connects the two variables using wire declarations. • Testbench: Here is a working testbench for a module that does the following: • Reads the input data from the control signals: module testbench(); input [3: 0] Data_Out; output [3: 0] Data_In; reg [3: 0] Data_In; reg MSB_In, LSB_In; // Get the input data from the control signals initial Data_In = 0; join initial begin fork join initial Data_In <= Data_Out[3]; join end fork join endmodule  This testbench uses wire declarations. It also uses reg variables. #### Testbenches that Verify initial reset The following test benches that verify the initial reset: module testbench(); reg rst; initial begin fork join fork join join end module  This testbenches does the following: • Assert the reset signal • De-assert the reset signal • Assert the reset signal • De-assert the reset signal The testbenches for the other test cases do the same thing. The module testbench() has a reg variable rst that is used to connect the reset signal to a control signal in the design. The following is the testbench: module testbench(); output [3: 0] Data_Out; reg [3: 0] Data_Out; initial fork begin initial Data_Out = 0; join initial Data_Out = 10'd12; join initial Data_Out = 0; join end module  This testbench does the following: • Assert the initial state • De-assert the state • Assert the initial state • De-assert the state The following testbench verifies the reset-on-the-fly: module testbench(); input [3: 0] Data_Out, Data_In; output [3: 0] Data_Out; initial fork begin initial Data_Out = 0; join initial Data_Out = 10'd12; join initial Data_Out = 0; join end module  This testbenches does the following: • Assert the initial state • De-assert the state • After 20ns, assert the state • De-assert