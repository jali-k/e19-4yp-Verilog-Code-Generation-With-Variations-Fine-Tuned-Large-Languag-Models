```verilog
module alu(s, A, B, F);
input [2:0] s;
input [3:0]