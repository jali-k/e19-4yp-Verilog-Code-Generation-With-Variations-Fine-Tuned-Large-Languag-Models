// Create a module containing a wire, reg, and assign statement
module reg_assign2( input in, output out );
    // Create the wire
    wire in1;
    // Create the registers
    reg output, reg_a;
    // Create the assign statement
    assign output = in1;
endmodule

### Verilog Code:
// Create a module containing a wire, reg, and assign statement
module reg_assign3