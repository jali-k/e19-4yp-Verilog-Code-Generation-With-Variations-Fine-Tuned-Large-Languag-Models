`module BubbleSort (input [3:0] data, output reg [3:0] data_sorted, output reg done);
always @* begin
    if (done