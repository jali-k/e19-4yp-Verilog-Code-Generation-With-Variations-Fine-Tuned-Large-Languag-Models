### Testbench File:
### Expected Output:

## How to Pack an Array of Packages:

To pack an array of packages, we apply the pack() function. It is used to pack an array. The pack() function is available in the package