module testbench ();
struct { bit[31:0] addr; } data;
always
begin
process
begin end
end
process data;
endmodule

### Variation Instruction:
Remove the always block and replace it with