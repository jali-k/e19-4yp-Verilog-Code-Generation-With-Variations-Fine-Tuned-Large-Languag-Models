### Verilog Code:
module muxdff(D0, D