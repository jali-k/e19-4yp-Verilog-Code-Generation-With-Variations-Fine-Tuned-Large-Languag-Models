always @(a[2:0]) begin
end
### Base Verilog Code:
always @(a[2:0]) begin  //$monitor triggers at t=0, t=2, t=5, t=6
end
`