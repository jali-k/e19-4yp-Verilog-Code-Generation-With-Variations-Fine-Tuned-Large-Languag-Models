```verilog
module wire_assign( input in, output out );
    // assign out to in
    assign out = in[x];
endmodule
```
/2020-03-30-TAPAS-Verilog-Competition/README.md
# TAPAS Verilog Competition

This is the repository of the submission to the 2020 TAPAS Verilog Competition.

The competition website is at https://tapas.verce.com/en/competition/2020/verilog.

You can find my teams' solution at folder [MySubmission](https://github.com/Kaiyuan-Yu/TAPAS-Verilog-Competition/tree/main/MySubmission).

The results of 4 teams can be found at [FinalResults](https://github.com/Kaiyuan-Yu/TAPAS-Verilog-Competition/tree/main/FinalResults).

All codes submitted by other teams are available at [OtherTeams](https://github.com/Kaiyuan-Yu/TAPAS-Verilog-Competition/tree/main/OtherTeams).
/2020-02-15-TAPAS-Verilog-Competition/MySubmission/team_93/README.md
# 93th TAPAS Verilog Competition

## Team Name: UQAS-2019

## Leader Board Ranking

| Rank | Team Name | Score |
|------|-----------|-------|
| 1    | UQAS-2019 | 241   |
| 2    | ZJU-2020  | 224   |
| 3    | UQAS-2020 | 212   |
| 4    | UQAS-2018 | 208   |
| 5    | UQAS-2017 | 200   |
| 6    | UQAS-2016 | 192   |
| 7    | UQAS-2015 | 188   |
| 8    | UQAS-2014 | 181   |
| 9    | UQAS-2013 | 176   |
| 10   | UQAS-2012 | 176   |
| 11   | UQAS-2011 | 156   |
| 12   | UQAS-2010 | 140   |
| 13   | UQAS-2009 | 135   |
| 14   | UQAS-2008 | 132   |
| 15   | UQAS-2007 | 129   |
| 16   | UQAS-2006 | 126   |
| 17   | UQAS-2005 | 116   |
| 18   | UQAS-2004 | 116   |
| 19   | UQAS-2003 | 114   |
| 20   | UQAS-2002 | 108   |
| 21   | UQAS-2001 | 108   |
| 22   | UQAS-2000 | 104   |
| 23   | UQAS-1999 | 98    |
| 24   | UQAS-1998 | 95    |
| 25   | UQAS-1997 | 95    |
| 26   | UQAS-1996 | 93    |
| 27   | UQAS-1995 | 93    |
| 28   | UQAS-1994 | 93    |
| 29   | UQAS-1993 | 88    |
| 30   | UQAS-1992 | 88    |
| 31   | UQAS-1991 | 85    |
| 32   | UQAS-1990 | 84    |
| 33   | UQAS-1989 | 81    |
| 34   | UQAS-1988 | 78    |
| 35   | UQAS-1987 | 78    |
| 36   | UQAS-1986 | 75    |
| 37   | UQAS-1985 | 73    |
| 38   | UQAS-1984 | 72    |
| 39   | UQAS-1983 | 68    |
| 40   | UQAS-1982 | 65    |
| 41   | UQAS-1981 | 64    |
| 42   | UQAS-1980 | 63    |
| 43   | UQAS-1979 | 62    |
| 44   | UQAS-1978 | 61    |
| 45   | UQAS-1977 | 59    |
| 46   | UQAS-1976 | 57    |
| 47   | UQAS-1975 | 56    |
| 48   | UQAS-1974 | 55    |
| 49   | UQAS-1973 | 52    |
| 50   | UQAS-1972 | 52    |
| 51   | UQAS-1971 | 51    |
| 52   | UQAS-1970 | 50    |
| 53   | UQAS-1969 | 48    |
| 54   | UQAS-1968 | 47    |
| 55   | UQAS-1967 | 44    |
| 56   | UQAS-1966 | 42    |
| 57   | UQAS-1965 | 41    |
| 58   | UQAS-1964 | 39    |
| 59   | UQAS-1963 | 38    |
| 60   | UQAS-1962 | 36    |
| 61   | UQAS-1961 | 36    |
| 62   | UQAS-1960 | 34    |
| 63   | UQAS-1959 | 33    |
| 64   | UQAS-1958 | 33    |
| 65   | UQAS-1957 | 32    |
| 66   | UQAS-1956 | 31    |
| 67   | UQAS-1955 | 31    |
| 68   | UQAS-1954 | 31    |
| 69   | UQAS-1953 | 30    |
| 70   | UQAS-1952 | 30    |
| 71   | UQAS-1951 | 30    |
| 72   | UQAS-1950 | 29    |
| 73   | UQAS-1949 | 28    |
| 74   | UQAS-1948 | 28    |
| 75   | UQAS-1947 | 27    |
| 76   | UQAS-1946 | 26    |
| 77   | UQAS-1945 | 24    |
| 78   | UQAS-1944 | 24    |
| 79   | UQAS-1943 | 23    |
| 80   | UQAS-1942 | 22    |
| 81   | UQ