module Clock_Prog(
input clk,
input [7:0] rstn
);

Clock_Prog M1 (clk, rstn);

endmodule