![Screen Shot 2022-11-02 at 09.31.52.png](data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABM0AAALRCAYAAAAkz1UaAAAMSGlDQ1BJQ0MgUHJvZmlsZQAASImVlwdUU1kagO97L73QAghICb0J0gkgJYQWQHoRbIQI2JFA7L3RAaTwAio8KqLgWgCxoqiIoGVlkEVCwLYs2KqiYkWx94UiCrp63nvn3jv3zXvfO/85c+bsmXPOwAJE9zwAoPeBudgUALjUy0tLBaAAkKADUk/GycsV5Ei4QgkWgPZT7/+XS5iLi/QaVz7nz/+/Sy+XcyEAAQiGQzgZArwMzg4BwB9FcqQKAJgL9Lt5LpKCAI1GZ7LZsP0CmEWKmBf4hbEaqL4DgJhMjGjmhQBgyBGgDwJAoACFgvz58c85/yU5ZYzM8Rjzj/8vx/zfUxY/wZs3MYwYs1HcDQC5iM941u3+f10j/y0xRwDgCQQZvJCJIKNBwjL5YhJHJhKQBQhgJ8YAIBLJyMxCfjYf4wY4Q2zh5wMHbAwgjg/wJTzBb2Ij3l4J2iZkdYGY7sOwDd0wz2JQeKIg7wzs2C9ykOwjP8Pz4zYjcYJRP5kQxhcCJQYJ4UHKHE6X+R/j4bL54xYZNlL2J8QhRgTq2Gnx/oL+M8UvWq134pIwWs3rRd9EfGSPy5Q/z+VyOqPWx6VxhW4XPFk/n9J2uHl+ZzpVKmGgxq+0nk7iM2qwkq5MnU97Q21/Tn5kDf5+fkN8gHrEZPwYNuoI2DgRYAJJwHu4uQZ59wHWyiXcw1zAB8IAEcgz4ALkQTfwA4p4NrT8ZDmBfB6CxRsYUeYEzGI8Bm4wDh9iP5K+znB16hmD/4gHp4iG4B9yIx89I7KZC+gVX023q8h/NxG0R+nOz1e48+4RX43wfqf+23vA/BKP+y3wR5h8JwM9kTjQQlhCCEGYI5rBfu+Oj5B70NtRCx4nXSbh+wGz5g81/N7/1PFhF4iC+F98Qq4fZm49Hh5v4t8t0A/yDQ716oF90I+21k4WTjJMtUm5f9/7H3nn9zFdWd/33dM2aWmSQhBZIlQEKH3jshCYTQQQMIImASM4iFYA4QyAQE4YAQEkI4QDgEwiEcAkmgY5jj7I/vXGfz3m9Xr1W7dnb3e5K+z36ec/Sj2lV1V63qWq26d2r5/aZtM1CmQOIJ8U3qc5HwNHFo4Ti+8ZL0x/ZY7nfqeO+K79hxw97Tv7Xn6fVd9z95nHnHqW9eVx377/l5XbWQ/fzD+L/9v/+3+qb1h3337Jz/3y+74Xn4/8388f/zf/x/Cj73+9/8/03+X8fu/3f//8f+x//3fR/50/3/9f/1/1v8//oF//9//P/3/+f/r/3f/P+P/8f+x/8f+h/+f5P/n+S/5//X/5//n/6//Z/8f+X/+//7//P/8/+r/2f+v/y//v/5//v/8//z/7P/7/1P8/2X8/8X/3/H/P+P/D/H/O/5//f/v/w//P//f9/9X/r/t/2f9//X/p/9P+f+X8f8P/r/u/wf/v+P/z/7/6f/3/z//v+P/u/7/7f/X/3/8//j/+f9v/3/7/7P8/3z/v+7/m/8f//8//x/9f/x//P8P/P8P/r/6/8f/B/8f/3//f/j//f8z/3/9/9n/P/3/Gf//5v8v/H/z/xv/v+H/5/+v/5/6/8H/H/7/wP/H/y/+f+X/j/9f/n/9/9n/P/z/yv/f/f8j/v/X/b/t/6f9/+v/F/6/+P/Z/z/5/+3/b/z/9P9n/v/w/y/8/+P/5/8X/3/2/+P/5/+v/z/7//n/5//3/X/7/5//3/f/1f9v/3/7//f/z/k/9P/D/6/9/8H/3/9/+f/V/x/+f/X/4f8P/n/x/5v/3/T/+//X/t/6f+z/2/8/+/8j/7/+/+n/d/+/6f+3/7/8/9//P/r/Hf9/8f83/L/7/5v/3/r/x/+v/z/7/xv/v+X/l/+//f+S/5/+f/f/4f/X/7/9/+P/L/8/+/3v8//T/+/+//H/1/+/+v/d/4/+f/f/r/7/+P/d/9/6f/L/2/+/+v/z/3/8/+z/X/3/7f/P/n/y/7P/H/6/8/+T/9/8/+T/t/8/+P/t/w/+f/H/8/8f/7/+//f/h/8//3/7/wf/v/n/t/w/8/+P/z/+f/n/5f9X/3/5/5H/f/j/1/+f/n/t/