module mux(sel, a, b, z);
parameter D = 1