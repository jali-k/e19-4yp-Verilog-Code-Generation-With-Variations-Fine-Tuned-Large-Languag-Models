module control_unit (flush_P0_P1, Ld_P1, Ld_P0, Ld, En, clock, rst);
output reg flush_P0_P1, Ld_P1, Ld_P0, Ld_R0;
input Ld, En, clock, rst;
reg [1: 0] state, next_state;
parameter S_idle = 0, S_1 = 1, S_full = 2, S_wait = 3;
always @ (posedge clock) if (rst) state <= S_idle;
else state <= next_state;
always @ (state, Ld, En) begin
flush_P0_P1 = 0;
Ld_P1 = 0;
Ld_P0 = 0;
Ld_R0 = 0;
next_state = S_idle;
case (state)
S_idle: if (En)
begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end
else flush_P0_P1 = 1;

S_1: begin next_state = S_full; Ld_P1 = 1; Ld_P0 = 1; end
S_full: if (Ld == 1) begin
Ld_R0 = 1;
case (En)
0: begin next_state = S_idle; flush_P0_P1 = 1; end
1: begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end
end
else begin
case (inside(x, state_table))
S_idle: next_state = S_idle;
S_1: next_state = S_1;
S_full: next_state = S_full;
S_wait: next_state = S_wait;
endcase
end
endcase
end
end

### Modified Top Level Code:
module top_level (clk, adata);
//...

clock clk;

//...

reg [31: 0] x;
reg [7: 0] y;
reg [1: 0] state, next_state;
reg En;
wire Ld, Rst;

//...

control_unit cu (En, Ld, Rst, clk, clk, state, next_state);
reg [1: 0] state, next_state;
reg En;
wire Ld, Rst;

//...

initial $display("state = %b, next_state = %b", state, next_state); x = 10010010010010010010010010010010; #10; // This code is repeated for each test case. while(1) begin #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; #10; clk = ~clk; end endmodule ### Hex-to-7seg Array Declaration: parameter [3: 0] state_table [7: 0] = {S_idle, S_1, S_full, S_wait, S_idle, S_1, S_full, S_wait}; ### Base Verilog Code: module control_unit (flush_P0_P1, Ld_P1, Ld_P0, Ld_R0, Ld, En, clock, rst); output reg flush_P0_P1, Ld_P1, Ld_P0, Ld_R0; input Ld, En, clock, rst; reg [1: 0] state, next_state; parameter S_idle = 0, S_1 = 1, S_full = 2, S_wait = 3; always @ (posedge clock) if (rst) state <= S_idle; else state <= next_state; always @ (state, Ld, En) begin flush_P0_P1 = 0; Ld_P1 = 0; Ld_P0 = 0; Ld_R0 = 0; next_state = S_idle; case (state) S_idle: if (En) begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end else flush_P0_P1 = 1; case (state) S_1: begin next_state = S_full; Ld_P1 = 1; Ld_P0 = 1; end S_full: if (Ld == 1) begin Ld_R0 = 1; case (En) 0: begin next_state = S_idle; flush_P0_P1 = 1; end 1: begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end end else next_state = S_wait; S_wait: if (Ld == 1) begin Ld_R0 = 1; case (En) 0: begin next_state = S_idle; flush_P0_P1 = 1; end 1: begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end end else next_state = S_wait; endcase endendmodule ### Variation Instruction: For the hex-to-7seg decoder, use `inside` to compare `x` against a constant array declared in dollar unit scope. ### Modified Code: module control_unit (flush_P0_P1, Ld_P1, Ld_P0, Ld_R0, Ld, En, clock, rst); output reg flush_P0_P1, Ld_P1, Ld_P0, Ld_R0; input Ld, En, clock, rst; reg [1: 0] state, next_state; parameter S_idle = 0, S_1 = 1, S_full = 2, S_wait = 3; always @ (posedge clock) if (rst) state <= S_idle; else state <= next_state; always @ (state, Ld, En) begin flush_P0_P1 = 0; Ld_P1 = 0; Ld_P0 = 0; Ld_R0 = 0; next_state = S_idle; case (state) S_idle: if (En) begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end else flush_P0_P1 = 1; case (state) S_1: begin next_state = S_full; Ld_P1 = 1; Ld_P0 = 1; end S_full: if (Ld == 1) begin Ld_R0 = 1; case (En) 0: begin next_state = S_idle; flush_P0_P1 = 1; end 1: begin next_state = S_1; Ld_P1 = 1; Ld_P0 = 1; end end else begin case (inside(x, state_table)) S_idle: next_state = S_idle; S_1: next_state = S_1; S_full: next_state = S_full; S_wait: next_state = S_wait; end end end endmodule ### Modified Top Level Code: module top_level (clk, adata); //... clock clk; //... //... reg [31: 0] x; reg [7: 0] y; reg [1: 0] state, next_state; reg En; wire Ld, Rst; //... control_unit cu (En, Ld, Rst, clk, clk, state, next_state); reg [1: 0] state, next_state; reg En; wire Ld, Rst; //... initial$display("state = %b, next_state = %b", state, next_state);
x = 10010010010010010010010010010010;
#10; // This code is repeated for each test case.
while(1) begin
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
#10;
clk = ~clk;
end
endmodule
### Hex-to-7