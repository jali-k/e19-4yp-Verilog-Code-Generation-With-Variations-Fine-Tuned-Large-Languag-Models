`decode_hex{16}` will compare x against 0.. 15.
`decode_hex{16: 0}` will compare x against 16.. 255.
`decode_hex{16: 16}` will compare x against 16.. 31.
`decode_hex{16: 16: 16}` will compare x against 16.. 31.
`decode_hex{8: 8}` will compare x against 8.. 15

## Lesson 7:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 7: Hex-to-7 Segment Decoder`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 8:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 8: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 9:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 9: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 10:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 10: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 11:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 11: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 12:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 12: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation/Projects/project1/Makefile
all:
	iverilog -D SIM -o testbench testbench.v
	vvp testbench
/Projects/project2/Makefile
all:
	iverilog -o testbench testbench.v
	vvp testbench

clean:
	rm -rf *.vcd
	rm -rf testbench
/Projects/project2/README.md
# Project 2 Code

##  and 

## Lesson 1:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 1: Hex-to-7 Segment Decoder`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 2:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 2: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 3:
1. Make sure to save your code in a.txt document
2. Make sure to save your code in a.zip file
2. Make sure to save your code in a.v file
3. Make sure you are modifying the code in a new Verilog file
4. Make sure to add the following to the top of your code:
`//  and 
// CE4507 - 001
// Lesson 3: Hex-to-7 Segment Decoder
// Purpose: Implement a hex-to-7 segment decoder and convert the hexadecimal 1A to the seven-segment representation in decimal 26`
### Simulation
1. Start your simulation
2. Wait for the simulation to finish
3. Click on the 'Results' icon in the top-right and select 'Save Waveform'
4. Save the file at a location that you choose
5. Close the simulation

## Lesson 4:
1. Make sure to save your code in a.txt document
2.