```verilog
typedef struct {
  rand bit [7:0] DataOut;
  bit [7:0] DataIn;
  bit ControlSignals;
} DataComponent;

module TestDataComponent(DataComponent_struct.DataOut, DataComponent_struct.DataIn, DataComponent_struct.ControlSignals);
DataComponent DataComponent_struct;
endmodule
```
In the "TestDataComponent" module, instead of `DataIn`, `DataOut`, and `ControlSignals`, you can now use the syntax `DataComponent_struct.DataOut`, `DataComponent_struct.DataIn`, `DataComponent_struct.ControlSignals`. Using this notation, we can access and modify the members of the struct.

Note: This will not generate any hardware. It's a structural Verilog design that uses a struct to represent the data component. Verilog also supports the use of classes for complex designs. However, the struct is a simpler construct and is typically used for simple, un-recursive data types.

Remember, the `rand` keyword in the struct will generate random values during the simulation, but you need to connect the struct to a testbench or another module to use it.

Also, keep in mind that using random variables should be used sparingly and not in critical paths of the design where a specific, repeatable sequence is required. This is primarily used for testbenches and simulations, not for actual hardware design. In hardware, the values of these variables usually come from the FPGA's fabric, not generated by the Verilog code.###

For example, you might have a testbench like this:

```verilog
module TestDataComponent (
  output [7:0] DataOut,
  input [7:0] DataIn,
  input ControlSignals
);

DataComponent DataComponent_struct;

initial begin
  #10; // Ensure the struct is ready
  $display("Random data output: %0d", DataComponent_struct.DataOut);
end

endmodule
```
In this example, the module will initialize the `DataOut` field of the struct with a random value, then print that value. This is often used for testing the randomization of the `DataOut` value.```