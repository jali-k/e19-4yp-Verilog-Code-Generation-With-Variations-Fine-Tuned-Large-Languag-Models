module netdelay1(x,y);
input x;
output [31:0] y; // output y as a unit width packed structure
wire #(2,1) [31:0] nn; // Declare wire 'nn' with rise=2, fall=1 delay
not (nn,x); // Assign NOT(x) to 'nn' (takes effect after rise/fall delay)
assign y=nn; // Assign 'nn' to 'y' (direct assignment)
endmodule
`

## Test Results

### Test Pass Result

All 6 Test Cases are Passed

### Test Case Result on Target Device

![](./images/test-result.png)

## Performance

### Target Device

#### Device Information

Verilog Model:

- Intel(R) FPGA Emulator for Windows with 128KB Cache and 256KB SRAM

#### Device Fmax Timing Constraints

![](./images/timing-const.png)

#### Device Fmax Timing Graph

![](./images/timing-graph.png)

#### Device Fmax Design Constraints

Fmax: 25.862001510946146

![](./images/design-const.png)

#### Device Fmax Design Graph

![](./images/design-graph.png)

### Compared with Other Solutions

All solutions can meet the constraints and design goals. However, we can observe some design details of the proposed design.

-  The proposed solution only needs 12 LUTs to realize the design of the network delay pipeline.
-  The proposed solution with 32 bit output bit width can achieve good timing while consuming only 16 LUTs.
-  The proposed solution with 32 bit output bit width can achieve good timing and design with 16 LUTs.

## Conclusion

Through this project, we have successfully constructed a network delay pipeline with Verilog and run the simulation on Intel FPGA Emulator. We have also analyzed the design details and compared with the existing design solutions. In this way, we can have more insights and knowledge on the design of the network delay pipeline on FPGA. We can also have more design inspiration.

## Reference

[Verilog HDL - Not Gate - W3SCHOOLS](https://www.w3schools.com/verilog/verilog_not.asp)

[How many LUTs does a NOT gate require?](https://electronics.stackexchange.com/questions/85795/how-many-luts-does-a-not-gate-require)

[HDL Design: A practical guide for beginner](https://ieeexplore.ieee.org/document/4012834)

[Verilog Tutorial](https://www.edaplayground.com/tutorials/verilog/verilog-tutorial-series-verilog-basics)

[Verilog Timing Constraints](https://www.allaboutcircuits.com/technical-articles/timing-constraints-in-verilog/)/Vivado/project/project.runs/impl_1/.vivado.mk
# Generated by Vivado on Thu Aug 19 14:37:14 CST 2021
# User: admin
# Date: 2021-08-19_14:37:27
# Flow: Sink
# Package: Vivado 2019.2
# IP Paint Size: 1080
# Command: C:/Program Files (x86)/Xilinx/Vivado/2019.2/bin/vivado -nojournal -nolog -mode batch -source..\..\netdelay1.tcl -tclargs

# Exit�Ą