module decoder4(A, B, AB, ABC, Q);
input