module tst_CMOSsw1();
	reg in,con; wire out;
	CMOSsw1 cmsw(out,in,con); // Instantiate CMOS switch
	initial begin in=1'b0; con=1'b1; end // Start enabled
	always #5 in =~in; // Toggle data
	always #3 con=~con; // Toggle control
	initial $monitor($time, "in = %b, con = %b, output = %b ",in,con,out);
	initial #20 $stop; // Stop simulation
endmodule
### Error Message:
$ ghdl -a tst_CMOSsw1.vhdl
tst_CMOSsw1.vhdl:24:16: warning: cannot determine value of expression:
  function result
    (in, con)
  end result
###