module SchedDelayA;
shortint a, b;
initial
begin
end
always @(b) a = b;
always @(a