### Base Code:
### Variation Instruction:
Modify the module definition and the assignment statements