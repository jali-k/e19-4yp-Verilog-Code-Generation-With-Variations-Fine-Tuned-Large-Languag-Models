module tst_CMOSsw1_1();
  reg in,con; wire out;
  CMOSsw1 cmsw(out,in,