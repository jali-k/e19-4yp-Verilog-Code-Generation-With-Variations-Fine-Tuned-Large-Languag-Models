module func4(x1, x2, x3, f);
input x