module top(output wire[7:0] s);
parameter n = 8;
wire[