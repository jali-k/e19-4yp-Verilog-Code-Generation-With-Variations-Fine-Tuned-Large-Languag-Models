- The two DFF will share the same clock.
  - Both DFF will toggle at the same time.
  - Both DFF will toggle at the same time even though they have different inputs.
  - The delay between the two DFF toggle can be seen in the waveform.
- ### Notes:
  - The two DFF will share the same clock.
  - Both DFF will toggle at the same time.
  - Both DFF will toggle at the same time even though they have different inputs.
  - The delay between the two DFF toggle can be seen in the waveform.