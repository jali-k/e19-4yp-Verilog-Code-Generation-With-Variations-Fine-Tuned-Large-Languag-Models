.
### Notes:
1.  The timing annotation is still correct.
2.  The code in the