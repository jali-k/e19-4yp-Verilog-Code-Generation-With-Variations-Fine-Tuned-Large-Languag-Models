```
always @(a, b, c, d, e, f, g, h) begin
...
end
```

## Test15: Xor9
### Description