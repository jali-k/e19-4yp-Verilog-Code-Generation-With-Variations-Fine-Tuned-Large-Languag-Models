module Problem1(input clk, di, output reg [3:0] sum);
  logic clk;
  logic di;
  always @(