module alu_6( output [3:0] d, output co,