module gates4_top (
input wire [3:0] sw,
output wire [2:0] ld
);
gates4 U1 (
.x(sw),
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0])
);
endmodule
module gates4_top (
input wire [3:0] sw,
output wire [2:0] ld
);
gates4 U1 (
.x(sw),
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0])
);
endmodule
module gates4_top (
input wire [3:0] sw,
output wire [2:0] ld
);
gates4 U1 (
.x(sw),
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0])
);
endmodule
module gates4_top (
input wire [3:0] sw,
output wire [2:0] ld
);
gates4 U1 (
.x(sw),
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0])
);
endmodule
module gates4_top (
input wire [3:0] sw,
output wire [2:0] ld
);
gates4 U1 (
.x(sw),
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0])
);
endmodule