module alu_tb (
input clk,
input alu,
input alu_op,
input [7:0] inA,
input [7:0] inB