module tst_nm_in();
  reg in; wire out;
  NMOSinv nmv(out,in); // Instantiate NMOS inverter
  initial
    in =1'b1; // Start with input high -> output low
  always
  initial $monitor($time, " in = %b, output = %b ",in,out);
  initial #15 $stop; // Stop simulation
endmodule
### Variation Description:
Add a case statement using inside with a function call used as an index into a 4D array.

The array consists of 24 sets of 3 rows of 8 NMOS inverters.  The array index is constructed using the functions from part 1 of this lab.  The "in" and "out" ports of the NMOSInverters are provided by the VHDL code as arguments to the NMOSInverter constructor.

The code reads 8 NMOS inverters at a time from the array and provides them with the input at the top of the array.  It then monitors the time and the values of the output ports of the inverters in the array.
### Test Output:
$ scoop -d 1 -l 128 -L 128 -L 64 -L 4 -L 2 -L 1  -f 1000  -m nm_in_out.txt nm_in_out.v
$ more nm_in_out.txt
# in  out
# --- ---
1000  1  0
1001  1  0
1002  1  0
1003  1  0
1004  1  0
1005  1  0
1006  1  0
1007  1  0
1008  1  0
1009  1  0
1010  1  0
1011  1  0
1012  1  0
1013  1  0
1014  1  0
1015  1  0
1016  1  0
1017  1  0
1018  1  0
1019  1  0
1020  1  0
1021  1  0
1022  1  0
1023  1  0
1024  1  0
1025  1  0
1026  1  0
1027  1  0
1028  1  0
1029  1  0
1030  1  0
1031  1  0
1032  1  0
1033  1  0
1034  1  0
1035  1  0
1036  1  0
1037  1  0
1038  1  0
1039  1  0
1040  1  0
1041  1  0
1042  1  0
1043  1  0
1044  1  0
1045  1  0
1046  1  0
1047  1  0
1048  1  0
1049  1  0
1050  1  0
1051  1  0
1052  1  0
1053  1  0
1054  1  0
1055  1  0
1056  1  0
1057  1  0
1058  1  0
1059  1  0
1060  1  0
1061  1  0
1062  1  0
1063  1  0
1064  1  0
1065  1  0
1066  1  0
1067  1  0
1068  1  0
1069  1  0
1070  1  0
1071  1  0
1072  1  0
1073  1  0
1074  1  0
1075  1  0
1076  1  0
1077  1  0
1078  1  0
1079  1  0
1080  1  0
1081  1  0
1082  1  0
1083  1  0
1084  1  0
1085  1  0
1086  1  0
1087  1  0
1088  1  0
1089  1  0
1090  1  0
1091  1  0
1092  1  0
1093  1  0
1094  1  0
1095  1  0
1096  1  0
1097  1  0
1098  1  0
1099  1  0
1100  1  0
1101  1  0
1102  1  0
1103  1  0
1104  1  0
1105  1  0
1106  1  0
1107  1  0
1108  1  0
1109  1  0
1110  1  0
1111  1  0
1112  1  0
1113  1  0
1114  1  0
1115  1  0
1116  1  0
1117  1  0
1118  1  0
1119  1  0
1120  1  0
1121  1  0
1122  1  0
1123  1  0
1124  1  0
1125  1  0
1126  1  0
1127  1  0
1128  1  0
1129  1  0
1130  1  0
1131  1  0
1132  1  0
1133  1  0
1134  1  0
1135  1  0
1136  1  0
1137  1  0
1138  1  0
1139  1  0
1140  1  0
1141  1  0
1142  1  0
1143  1  0
1144  1  0
1145  1  0
1146  1  0
1147  1  0
1148  1  0
1149  1  0
1150  1  0
1151  1  0
1152  1  0
1153  1  0
1154  1  0
1155  1  0
1156  1  0
1157  1  0
1158  1  0
1159  1  0
1160  1  0
1161  1  0
1162  1  0
1163  1  0
1164  1  0
1165  1  0
1166  1  0
1167  1  0
1168  1  0
1169  1  0
1170  1  0
1171  1  0
1172  1  0
1173  1  0
1174  1  0
1175  1  0
1176  1  0
1177  1  0
1178  1  0
1179  1  0
1180  1  0
1181  1  0
1182  1  0
1183  1  0
1184  1  0
1185  1  0
1186  1  0
1187  1  0
1188  1  0
1189  1  0
1190  1