<img src="https://raw.githubusercontent.com/ShubhamGupta01/Randomization/master/img/proc.PNG" alt="Randomization" width="500">
### Results:
<img src="https://raw.githubusercontent.com/ShubhamGupta01/Randomization/master/img/proc%20Result.PNG" alt="Results" width="500">### Base Verilog Code:
module testbench ();
generate data;
process data;
endmodule
### Variation Instruction:
Replace the data construct with an alternativ