module show_aa(ao,ai);
  output logic ao;
  input show_aa_aa_t ai;
  wire logic ao;
  show_aa_aa_t ao;
  wire logic ai;
  show_aa_aa_t ai;
  not #2 (ao,ai);
endmodule