module tst_wand1; //testbench
reg i1,i2;
wire o;
wand1 ww(i1,i2,o);
wire [3:0] tmp; // added tmp
initial
begin
i1=0; i2=0;
tmp=~i1; // Drv1=pull0, Drv2=pull0 -> o = pull0 (wand rule)
end
initial $monitor($time,"i1=%b,i2=%b,o=%b",i1,i2,tmp[1:0]); // Changed to tmp[1:0]
initial $stop;
endmodule

And the output:

i1=0000 i2=0000 o=00
i1=0000 i2=0001 o=01
i1=0000 i2=0010 o=10
i1=0000 i2=0011 o=11
i1=0000 i2=0100 o=10
i1=0000 i2=0101 o=11
i1=0000 i2=0110 o=11
i1=0000 i2=0111 o=11
i1=0000 i2=1000 o=00
i1=0000 i2=1001 o=01
i1=0000 i2=1010 o=01
i1=0000 i2=1011 o=01
i1=0000 i2=1100 o=01
i1=0000 i2=1101 o=01
i1=0000 i2=1110 o=01
i1=0000 i2=1111 o=01
i1=0001 i2=0000 o=00
i1=0001 i2=0001 o=00
i1=0001 i2=0010 o=00
i1=0001 i2=0011 o=01
i1=0001 i2=0100 o=10
i1=0001 i2=0101 o=11
i1=0001 i2=0110 o=11
i1=0001 i2=0111 o=11
i1=0001 i2=1000 o=10
i1=0001 i2=1001 o=11
i1=0001 i2=1010 o=11
i1=0001 i2=1011 o=11
i1=0001 i2=1100 o=11
i1=0001 i2=1101 o=11
i1=0001 i2=1110 o=11
i1=0001 i2=1111 o=11
i1=0010 i2=0000 o=00
i1=0010 i2=0001 o=00
i1=0010 i2=0010 o=00
i1=0010 i2=0011 o=01
i1=0010 i2=0100 o=10
i1=0010 i2=0101 o=11
i1=0010 i2=0110 o=11
i1=0010 i2=0111 o=11
i1=0010 i2=1000 o=10
i1=0010 i2=1001 o=11
i1=0010 i2=1010 o=11
i1=0010 i2=1011 o=11
i1=0010 i2=1100 o=11
i1=0010 i2=1101 o=11
i1=0010 i2=1110 o=11
i1=0010 i2=1111 o=11
i1=0011 i2=0000 o=00
i1=0011 i2=0001 o=00
i1=0011 i2=0010 o=00
i1=0011 i2=0011 o=01
i1=0011 i2=0100 o=10
i1=0011 i2=0101 o=11
i1=0011 i2=0110 o=11
i1=0011 i2=0111 o=11
i1=0011 i2=1000 o=10
i1=0011 i2=1001 o=11
i1=0011 i2=1010 o=11
i1=0011 i2=1011 o=11
i1=0011 i2=1100 o=11
i1=0011 i2=1101 o=11
i1=0011 i2=1110 o=11
i1=0011 i2=1111 o=11
i1=0100 i2=0000 o=00
i1=0100 i2=0001 o=00
i1=0100 i2=0010 o=00
i1=0100 i2=0011 o=01
i1=0100 i2=0100 o=10
i1=0100 i2=0101 o=11
i1=0100 i2=0110 o=11
i1=0100 i2=0111 o=11
i1=0100 i2=1000 o=10
i1=0100 i2=1001 o=11
i1=0100 i2=1010 o=11
i1=0100 i2=1011 o=11
i1=0100 i2=1100 o=11
i1=0100 i2=1101 o=11
i1=0100 i2=1110 o=11
i1=0100 i2=1111 o=11
i1=0101 i2=0000 o=00
i1=0101 i2=0001 o=00
i1=0101 i2=0010 o=00
i1=0101 i2=0011 o=01
i1=0101 i2=0100 o=10
i1=0101 i2=0101 o=11
i1=0101 i2=0110 o=11
i1=0101 i2=0111 o=11
i1=0101 i2=1000 o=10
i1=0101 i2=1001 o=11
i1=0101 i2=1010 o=11
i1=0101 i2=1011 o=11
i1=0101 i2=1100 o=11
i1=0101 i2=1101 o=11
i1=0101 i2=1110 o=11
i1=0101 i2=1111 o=11
i1=0110 i2=0000 o=00
i1=0110 i2=0001 o=00
i1=0110 i2=0010 o=00
i1=0110 i2=0011