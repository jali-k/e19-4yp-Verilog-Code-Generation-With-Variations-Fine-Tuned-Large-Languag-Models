module IR ( input [7:0] data_in, input load, clk,
output reg [7:0] data_out );
// Simple register (Instruction Register) loaded on posedge clk when load is high
always @( posedge clk )
if ( load ) data_out <= data_in; // 1D array
data_out <= data_in; // 2D array
data_out <= data_in[1]; // 3D array
data_out <= data_in[1:3]; // 4D array
endmodule
To test the variations, modify the top-level testbench module as follows:
module tb_IR ( );
... // Other testbench code...
reg [7:0] data_in;
reg load;
reg clk;
assign clk = 1'b0;
generate
// Single-Dimensional array (one-dimensional logic-vector)
for ( data_in = 0; data_in <= 255; data_in++ )
begin
assign data_in = data_in;
assign clk = 0;
assign load = 1;
// 2D array (two-dimensional logic-vector)
for ( data_in = 0; data_in <= 511; data_in += 32 )
begin
assign data_in = data_in;
assign clk = 0;
assign load = 1;
// 3D array (three-dimensional logic-vector)
for ( data_in = 0; data_in <= 1023; data_in += 1024 )
begin
assign data_in = data_in;
assign clk = 0;
assign load = 1;
// 4D array (four-dimensional logic-vector)
for ( data_in = 0; data_in <= 2047; data_in += 2048 )
begin
assign data_in = data_in;
assign clk = 0;
assign load = 1;
end
end
assign clk = 1;
assign load = 0;
end
end
endmodule
After running the testbench, use waveform viewer to verify the generated waveforms as follows:
141
142
143
144
145
146
147
148
149
150
151
152
153
154
155
156
157
158
159
160
161
162
163
164
165
166
167
168
169
170
171
172
173
174
175
176
177
178
179
180
181
182
183
184
185
186
187
188
189
190
191
192
193
194
195
196
197
198
199
200
201
202
203
204
205
206
207
208
209
210
211
212
213
214
215
216
217
218
219
220
221
222
223
224
225
226
227
228
229
230
231
232
233
234
235
236
237
238
239
240
241
242
243
244
245
246
247
248
249
250
251
252
253
254
255
256
257
258
259
260
261
262
263
264
265
266
267
268
269
270
271
272
273
274
275
276
277
278
279
280
281
282
283
284
285
286
287
288
289
290
291
292
293
294
295
296
297
298
299
300
301
302
303
304
305
306
307
2018  and 
308
...
318
319
320
321
322
323
324
325
326
327
328
329
330
331
332
333
334
335
336
337
338
339
340
341
342
343
344
345
346
347
348
349
350
351
352
353
354
355
356
357
358
359
360
361
362
363
364
365
366
367
368
369
370
371
372
373
374
375
376
377
378
379
380
381
382
383
384
385
386
387
388
389
390
391
392
393
394
395
396
397
398
399
400
401
402
403
404
405
411
412
413
414
415
416
417
418
419
520
421
422
423
424
425
426
427
428
429
430
431
432
433
434
435
436
437
438
439
440
441
442
443
444
445
446
447
448
449
450
451
452
453
454
455
456
457
458
459
460
461
462
463
464
465
466
467
468
469
470
471
472
473
474
475
476
477
478
479
480
481
482
483
484
485
486
487
488
489
490
491
492
493
494
495
496
497
498
499
500
501
502
503
504
505
506
507
508
509
510
511
512
513
514
515
516
517
518
519
520
521
522
523
524
525
526
527
528
529
530
531
532
533
534
535
536
53