```
// Check XMR usage
if(BCD_in inside { pkg