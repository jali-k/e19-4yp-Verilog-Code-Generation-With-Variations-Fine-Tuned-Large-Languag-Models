// Create a module with one input and one output that behaves like a reg
module logic_assign(