#### Include Solution: