module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module ALU2 (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
module MyModule (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
specify
    specify
    specify
    specparam tRise = 5, tFall = 4;
    (Clk *> Result) = (tRise, tFall);
    (Clk *> ArgA) = (tRise, tFall);
    (Clk *> ArgB) = (tRise, tFall);
    (Clk *> ArgA) = (tRise, tFall);
    (Clk *> ArgB) = (tRise, tFall);
    (Clk *> ArgA) = (tRise, tFall);
    (Clk *> ArgB) = (tRise, tFall);
    (Clk *> ArgA) = (tRise, tFall);
    (Clk *> ArgB) = (tRise, tFall);
    (Clk *> ArgA) = (tRise, tFall);