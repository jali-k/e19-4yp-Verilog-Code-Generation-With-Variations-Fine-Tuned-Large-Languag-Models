```
module