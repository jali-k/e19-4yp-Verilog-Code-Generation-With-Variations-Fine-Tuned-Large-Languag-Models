module latch (input d, c, output q, q_b );
input [7:0] d;
input c;
output reg [7