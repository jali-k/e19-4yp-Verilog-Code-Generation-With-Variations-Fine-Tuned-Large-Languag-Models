module dff(do,di,