module t_decoder();
input a, b, c;
wire [4:0] d;
wire [4:0] d0, d1, d2, d