module wire_assign( input bit in, output out );
    assign out = in;
endmodule
### Results:
The output is a 1-bit (bit) with the same value as the input in