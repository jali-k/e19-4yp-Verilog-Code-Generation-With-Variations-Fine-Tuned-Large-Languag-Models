module wire_assign( input bit in, output bit out );
    // assign out to in
    assign out = in;
endmodule