module Problem9(input [3:0] a, b, output [3:0] sum);
  reg x = 4'b0110, y = 4'b01