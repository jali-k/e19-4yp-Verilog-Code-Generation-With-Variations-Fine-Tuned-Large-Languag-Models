module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;// a1,a2,b1,b2 form the input
//ports of the module
output o;//o is the single output port of the module
wire o1,o2;//o1 and o2 are intermediate signals
//within the module
and g1(o1,a1,a2); //The AND gate primitive has two
and g2(o2,b1,b2);// instantiations with assigned
//names g1 & g2.
nor g3(o,o1,o2);//The nor gate has one instantiation
//with assigned name g3.
endmodule
### SMT-LIB-v2:
(assert (or  a1 a2 b1 b2 (and a2 b1 b2)))
(assert (or  a1 a2 b1 b2 (and a1 b2 b1)))
(assert (or  a1 a2 b1 b2 (and a2 b2 a1)))
(assert (or  a1 a2 b1 b2 (and a1 b1 a2)))
(assert (or  a1 a2 b1 b2 (and a1 b1 a2)))
(assert (or  a1 a2 b1 b2 (and a1 b1 b2)))
(assert (or  a1 a2 b1 b2 (and a1 a2 b1)))
(assert (or  a1 a2 b1 b2 (and a2 a1 b1)))
(assert (or  a1 a2 b1 b2 (and a2 a1 b2)))
(assert (or  a1 a2 b1 b2 (and a1 a2 a1)))
(assert (or  a1 a2 b1 b2 (and a1 a2 a2)))
(assert (or  a1 a2 b1 b2 (and a1 b1 b1)))
(assert (or  a1 a2 b1 b2 (and a1 b1 b2)))
(assert (or  a1 a2 b1 b2 (and a1 b2 b1)))
(assert (or  a1 a2 b1 b2 (and a2 b1 b1)))
(assert (or  a1 a2 b1 b2 (and a2 b1 b2)))
(assert (or  a1 a2 b1 b2 (and a2 b2 b1)))
(assert (or  a1 a2 b1 b2 (and b1 b1 b1)))
(assert (or  a1 a2 b1 b2 (and b1 b1 b2)))
(assert (or  a1 a2 b1 b2 (and b1 b2 b1)))
(assert (or  a1 a2 b1 b2 (and b2 b1 b1)))
(assert (or  a1 a2 b1 b2 (and b2 b1 b2)))
(assert (or  a1 a2 b1 b2 (and b2 b2 b1)))
(assert (or  a1 a2 b1 b2 (and b2 b2 b2)))
(check-sat)
(get-model)
### Veri-fu result:
This Veri-fu run is successful
### SMT-LIB-v2:
(assert (and  a1 a1 a1))
(assert (and  a1 a1 a2))
(assert (and  a1 a2 a1))
(assert (and  a1 a2 a2))
(assert (and  a1 a2 b1))
(assert (and  a1 a2 b2))
(assert (and  a1 a2 b1))
(assert (and  a1 a2 b2))
(assert (and  a1 b1 b1))
(assert (and  a1 b1 b2))
(assert (and  a1 b2 b1))
(assert (and  a1 b2 b2))
(assert (and  a2 b1 b1))
(assert (and  a2 b1 b2))
(assert (and  a2 b2 b1))
(assert (and  a2 b2 b2))
(check-sat)
(get-model)
### Veri-fu result:
This Veri-fu run is successful
### SMT-LIB-v2:
(assert (= a0 (and b1 b2)))
(assert (= a2 (and a1 b2)))
(assert (= a1 (and a2 b1)))
(assert (= a1 (and a2 b2)))
(assert (= a2 (and a1 b1)))
(assert (= a1 (and a1 b1)))
(assert (= a1 (and a1 b2)))
(assert (= a0 (and a1 b1)))
(assert (= a0 (and a2 b1)))
(assert (= a1 (and a2 b2)))
(assert (= a0 (and a1 a1)))
(assert (= a2 (and a1 a2)))
(assert (= a0 (and a2 a1)))
(assert (= a1 (and a2 a2)))
(assert (= a2 (and a1 b2)))
(assert (= a2 (and a2 b2)))
(assert (= a0 (and a2 b2)))
(assert (= a1 (and a1 b1)))
(assert (= a2 (and a1 b2)))
(assert (= a0 (and a1 b2)))
(assert (= a0 (and a2 b1)))
(assert (= a0 (and a2 b2)))
(assert (= a1 (and a2 b1)))
(assert (= a1 (and a2 b2)))
(assert (= a0 (and a2 b1)))
(assert (= a0 (and a1 b1)))
(assert (= a1 (and a1 b2)))
(assert (= a2 (and a2 b2)))
(assert (= a1 (and a1 b1)))
(assert (= a2 (and a1 b1)))
(assert (= a1 (and a1 b2)))
(assert (= a2 (and a2 b1)))
(assert (= a2 (and a2 b2)))
(assert (= a2 (and a1 a2)))
(assert (= a0 (and a1 a2)))
(assert (= a0 (and a2 a1)))
(assert (= a0 (and a2 a2)))
(assert (= a1 (and a1 a1)))
(assert (= a0 (and a1 a1)))
(assert (= a2 (and a1 a2)))
(assert (= a1 (and a1 a2)))
(assert (= a0 (and a1 a1)))
(assert (= a2 (and a2 a1)))
(assert (= a2 (and a2 a2)))
(assert (> (and a1 b1 b1) a0))
(assert (> (and a1 b1 b2) a0))
(assert (> (and a1 b2 b1) a0))
(assert (> (and a1 b2 b2) a0))
(assert (> (and a2 b1 b1) a0))
(assert (> (and a2 b1 b2) a0))
(assert (> (and a2 b2 b1) a0))
(assert (> (and a2 b2 b2) a0))
(assert (> (and a1 a1 b1) a0))
(assert (> (and a1 a1 b2) a0))
(assert (> (and a1 b1 b1) a0))
(assert (> (and a1 b1 b2) a0))
(assert (> (and a1 b2 b1) a0))
(assert (> (and a1 b2 b2) a0))
(assert (> (and a2 b1 b1) a0))
(assert (> (and a2 b1 b2) a0))
(assert (> (and a2 b2 b1) a0))
(assert (> (and a2 b2 b2) a0))
(assert (> (and a1 b1 a1) a0))
(assert (> (and a1 b1 a2) a0))
(assert (> (and a1 a2 b1) a0))
(assert (> (and a1 a2 b2) a0))
(assert (> (and a1 a2 a1) a0))
(assert (> (and a1 a2 a2) a0))
(assert (> (and b1 b1 b1) a0))
(assert (> (and b1 b1 b2) a0))
(assert (> (and b1 b2 b1) a0))
(assert (> (and b1 b2 b2) a0))
(assert (> (and b2 b1 b1) a