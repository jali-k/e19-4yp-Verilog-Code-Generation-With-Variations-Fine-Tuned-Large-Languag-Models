module Anding (input a, b, output y);
and (y, a, b);
endmodule
### Expected Output:
```
module Anding (input a, b, output y);
and (y, a, b);
endmodule
```

### Score: 100
### Test Cases Passed: 3