reg_array[2] = reg_array[2] | reg_array2[0];

### Expected Output: