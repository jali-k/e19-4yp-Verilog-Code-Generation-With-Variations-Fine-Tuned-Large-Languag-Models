// Verilog code for Problems 5
// modified to use a