module tb_sw2led2;

reg [7:0] sw;
wire [7:0] ld;

signed_led2 led2(.sw(sw),.ld(ld));

initial begin
    sw = 0;
    #100;
    sw = 8'b00000001;
    #100;
    sw = 8'b00000010;
    #100;
    sw = 8'b00000011;
    #100;
    sw = 8'b00000100;
    #100;
    sw = 8'b00000101;
    #100;
    sw = 8'b00000110;
    #100;
    sw = 8'b00000111;
    #100;
    sw = 8'b00001000;
    #100;
    sw = 8'b00001001;
    #100;
    sw = 8'b00001010;
    #100;
    sw = 8'b00001011;
    #100;
    sw = 8'b00001100;
    #100;
    sw = 8'b00001101;
    #100;
    sw = 8'b00001110;
    #100;
    sw = 8'b00001111;
    #100;
    sw = 8'b00010000;
    #100;
    sw = 8'b00010001;
    #100;
    sw = 8'b00010010;
    #100;
    sw = 8'b00010011;
    #100;
    sw = 8'b000