```
module nil;
reg [3:0] a