```verilog
module show_aa(
    ao, ai, bi, bo
); 

    output a