module dec2_4beh(q,i);
output [3:0] q;
input [1:0]i;