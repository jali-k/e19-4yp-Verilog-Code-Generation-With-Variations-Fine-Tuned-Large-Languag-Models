class schedDelayA_t #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends $clog2(MAX_INPUT); endclass reg [MAX_INPUT-1:0]a; wire [MAX_OUTPUT-1:0]a_; reg [MAX_INPUT-1:0]b; wire [MAX_OUTPUT-1:0]b_; initial begin for (genvar i=0; i<MAX_INPUT; i=$clog2(MAX_INPUT)-1; i>=0)
begin
end
for (genvar i=0; i<MAX_INPUT; i=$clog2(MAX_INPUT)-1; i>=0) begin a[i] = i==1'b1? 1'bx : 1'b0; b[i] = i==1'b1? 1'b1 : 1'bx; end for (genvar i=0; i<MAX_OUTPUT; i=$clog2(MAX_OUTPUT)-1; i>=0)
begin
end
for (genvar i=0; i<MAX_OUTPUT; i=$clog2(MAX_OUTPUT)-1; i>=0) begin assign a_ = a[i]; assign b_ = b[i]; end for (genvar i=0; i<MAX_OUTPUT; i=$clog2(MAX_OUTPUT)-1; i>=0)
begin
end
endmodule

class schedDelayA_t_inst0 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_test #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst1 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst2 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst3 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst4 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst5 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst6 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst7 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst8 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst9 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst10 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst11 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst12 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst13 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst14 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst15 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst16 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst17 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst18 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst19 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst20 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst21 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst22 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst23 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst24 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst25 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst26 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst27 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst28 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst29 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst30 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst31 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst32 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t #(MAX_INPUT, MAX_OUTPUT);
endclass

class schedDelayA_t_inst33 #(parameter int MAX_INPUT = 5, parameter int MAX_OUTPUT = 5)
extends schedDelayA_t