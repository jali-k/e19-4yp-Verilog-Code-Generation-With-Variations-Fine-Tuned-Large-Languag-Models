module mixed_sim;
reg dcontrol, x, y;
reg [31:0] data;
reg [31:0] bus;