module reg4(Sum, Clock, Reset, RegSum);
input [3:0] RegSum;
input Clock, Reset;
output [3:0] Sum;
wire [3:0] Sum;
reg [3:0