```
`inside {S_4, S_8}
```