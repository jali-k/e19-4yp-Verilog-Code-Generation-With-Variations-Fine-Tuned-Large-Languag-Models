module tst_ctr_wt;
reg clk;
assign clk=clk+1;
reg[3:0]N;
wire[3:0]a;

`assign N=inside(a,0,10,1);`

`assign N=inside(a,5,7,1);`

`assign N=inside(a,0,10,2);`

`assign N=inside(a,0,10,4);`

`assign N=inside(a,0,10,7);`

`assign N=inside(a,0,10,8);`

`assign N=inside(a,0,10,10);`

`assign N=inside(a,0,3,1);`

`assign N=inside(a,3,5,1);`

`assign N=inside(a,1,3,1);`

`assign N=inside(a,3,3,1);`

`assign N=inside(a,0,3,2);`

`assign N=inside(a,3,3,2);`

`assign N=inside(a,2,2,2);`

`assign N=inside(a,5,7,2);`

`assign N=inside(a,2,2,4);`

`assign N=inside(a,1,1,4);`

`assign N=inside(a,9,9,4);`

`assign N=inside(a,5,7,7);`

`assign N=inside(a,8,8,7);`

`assign N=inside(a,5,5,7);`

`assign N=inside(a,8,8,8);`

`assign N=inside(a,1,1,8);`

`assign N=inside(a,9,9,8);`

`assign N=inside(a,5,5,8);`

`assign N=inside(a,0,9,2);`

`assign N=inside(a,0,9,4);`

`assign N=inside(a,0,9,7);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=inside(a,9,2,10);`

`assign N=inside(a,9,1,10);`

`assign N=inside(a,0,8,10);`

`assign N=inside(a,0,2,10);`

`assign N=inside(a,0,1,10);`

`assign N=inside(a,1,10,10);`

`assign N=inside(a,9,9,10);`

`assign N=inside(a,9,4,10);`

`assign N=inside(a,9,3,10);`

`assign N=