```
class FSM;
    parameter bool A = 0, B = 1;
    parameter uint FSM_STATE_COUNT;
    parameter FSM_STATE_COUNT;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] FSM_STATE_TYPE;
    typedef logic [FSM_STATE_COUNT-1:0] F