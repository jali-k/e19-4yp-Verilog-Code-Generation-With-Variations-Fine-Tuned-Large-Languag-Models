// Verilog Code:
module show_aa(ai); // NOT gate with delay 2
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  //output ao; input ai; pack packed ai;
  output ao; input ai; pack packed ai;
  not #2 (ao,ai);
endmodule
// Java Code:
class show_aa {
    int ao;
    //int ai;