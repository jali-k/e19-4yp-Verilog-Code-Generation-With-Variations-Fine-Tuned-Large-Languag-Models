module par(in, parity, all_ones);
input [