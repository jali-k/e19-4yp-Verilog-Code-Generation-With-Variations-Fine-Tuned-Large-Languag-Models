module and2(a, b, f);
input a, b;
output signed f;
assign f = a & b;
endmodule

## Question 11:
Implement the following circuit using the four-input CMOS NAND gate described in the Karnaugh map below:

![Q11](https://github.com/babyvibes/ECE6122/blob/7f9d9a4fddb8c99831df60947715