### Test Vector:
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
32'h890abcde  32'h1234abcd  32'h33333333  32'h890abcde
#### Simulation Results:
Test Number 0:
The first test case is for unsigned addition.
A = 32'h890abcde, B = 32'h1234abcd, result = 32'h9b3ebce6, carry = 0, zero = 0
The test passed!

Test Number 1:
The second test case is for unsigned subtraction.
A = 32'h1234abcd, B = 32'h890abcde, result = 32'he6d85031, carry = 0, zero = 0
The test passed!

Test Number 2:
The third test case is for unsigned multiplication.
A = 32'h1234abcd, B = 32'h890abcde,