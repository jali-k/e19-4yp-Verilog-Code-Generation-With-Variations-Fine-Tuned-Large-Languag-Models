`timescale 1ns/100ps
module ALU8 (input [7:0] left, right, input [1:0] mode, output reg [7:0] ALUout);
always_comb begin
    ALUout = {left[7], left[6:0], left[5], left[3:0], left[2], left[1:0]};
    case (mode)
        0: ALUout = [left[7], left[6:0], left[5], left[3:0], left[2], left[1:0]] + [right[7], right[6:0], right[5], right[3:0], right[2], right[1:0]];
        1: ALUout = [left[7], left[6:0], left[5], left[3:0], left[2], left[1:0]] - [right[7], right[6:0], right[5], right[3:0], right[2], right[1:0]];
        2: ALUout = [left[7], left[6:0], left[5], left[3:0], left[2], left[1:0]] & [right[7], right[6:0], right[5], right[3:0], right[2], right[1:0]];
        3: ALUout = [left[7], left[6:0], left[5], left[3:0], left[2], left[1:0]] | [right[7], right[6:0], right[5], right[3:0], right[2], right[1:0]];
        default: ALUout = 8'bx;
    endcase
end

endmodule
### Execution:
```
% vcs dut.v
%./simv 
% run 1000000
% vvp -modname dut -full64 simv.vcd | grep ALUout
ALUout=d008
ALUout=d008
ALUout=d000
ALUout=d008
ALUout=d008
ALUout=d000
ALUout=d008
ALUout=d000
ALUout=d000
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d000
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d000
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d000
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d000
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d008
ALUout=d00