module IR_tb( );
localparam NUM_BITS = 7;
localparam NUM_BYTES = 8;

// Input 
reg [NUM