module Fibonacci_gen;
reg [15:0] Fibonacci;
reg [15:0] F_1;
reg [15:0] F_2;
reg [15:0] index;
reg [7:0] F_index;
reg [7:0] F_1_index;
reg [7:0] F_2_index;
wire [7:0] index_reg;
wire [7:0