module Oring (myunion);
	input [1:0] a, b;
	output y;
	wire [1:0] out_myuniona;
	wire [1:0] out_myunionb;
	wire [1:0] out_y;
	Anding #(.y(out_myuniona)) myanding_a(.a(a[1]),.b(a[0]));
	Anding #(.y(out_myunionb)) myanding_b(.a(b[1]),.b(b[0]));
	Oring #(.y(out_y)) myor(.a(out_myuniona),.b(out_myunionb));
	assign y = out_y;
endmodule
### New Input Signal:
```
myunion:  {
	a: {
		type: "input",
		name: "a",
		value: "0",
		width: 2,
		base: "DEC"
	},
	b: {
		type: "input",
		name: "b",
		value: "0",
		width: 2,
		base: "DEC"
	},
}
```
### Expected Output:
```
% iverilog -o test.vvp myunion.v test.v
% vvp test.vvp
% vvp -M. -m iverilog_testsuite myunion.v test.v
%
% 0
% 1
% 2
% 3
% 4
```
### Expected Testbench Code:
```
initial begin
	$dumpfile("myunion.vpd");
	$dumpvars(0, myunion);
	#1 a = "0";
	#1 a = "1";
	#1 a = "2";
	#1 a = "3";
	#1 a = "4";
	$finish;
end
```
### Generated Verilog:
```
module myunion (a, b, y);
	input [1:0] a;
	input [1:0] b;
	output [1:0] y;
	Anding myanding_a (.a(a[1]),.b(a[0]),.y(myunion_a));
	Anding myanding_b (.a(b[1]),.b(b[0]),.y(myunion_b));
	Oring myor (.a(myunion_a),.b(myunion_b),.y(y));
endmodule
```
### Verilator Generated Testbench:
```
#include <verilated.h>
#include "Vmyunion.h"

int
main()
{
    Verilated::commandArgs(1, "myunion.v");
    Vmyunion* tb = new Vmyunion;

    // Initialize Verilator variables
    tb->a = 0;
    tb->b = 0;

    // Tick clock until simulation is finished
    int clock = 0;
    while (!Verilated::gotFinish()) {
        tb->eval();

        // Dump the testbench state to a vcd file
        tb->trace(VCD_C::vcdPopt(Verilated::traceEver()));
        tb->trace(VCD_C::vcdPopt(Verilated::traceEver()));
        tb->trace(VCD_C::vcdPopt(Verilated::traceEver()));
        tb->trace(VCD_C::vcdPopt(Verilated::traceEver()));
        tb->trace(VCD_C::vcdPopt(Verilated::traceEver()));

        // Increment clock by one
        clock++;
    }

    // Close the trace
    tb->trace(NULL, 0);

    // Clean up the simulation
    delete tb;
    exit(0);
}
```
### Expected Test Vectors:
```
% iverilog -o test.vvp myunion.v test.v
% vvp test.vvp
% vvp -M. -m iverilog_testsuite myunion.v test.v
%
% 0
% 1
% 2
% 3
% 4
```
### Test Vectors Generated by Icarus Verilog:
```
.input a
.input b
.output y

#1 a = "0";
#1 a = "1";
#1 a = "2";
#1 a = "3";
#1 a = "4";
```
/lib/src/verilog/printer/VerilogPrinter.h
//
// Copyright (C) [2020] Futurewei Technologies, Inc.
//
// FORCE-RISCV is licensed under the Apache License, Version 2.0 (the "License");
//  you may not use this file except in compliance with the License.
//  You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
// THIS SOFTWARE IS PROVIDED ON AN "AS IS" BASIS, WITHOUT WARRANTIES OF ANY KIND, EITHER
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO NON-INFRINGEMENT, MERCHANTABILITY OR
// FIT FOR A PARTICULAR PURPOSE.
// See the License for the specific language governing permissions and
// limitations under the License.
//
#ifndef _VERILOG_PRINTER_H
#define _VERILOG_PRINTER_H

#include <ostream>

#include "GenPrinter.h"
#include "Object.h"

namespace Force {

  class AIG;
  class AIGNode;
  class AIGNodeSet;
  class AIGVector;
  class AIGVectorSet;
  class AIGVariableNode;
  class AIGVariableNodeSet;
  class AIGVariableVector;
  class AIGVariableVectorSet;
  class BitVector;
  class BitVectorSet;
  class CodeNode;
  class CodeNodeSet;
  class Constraint;
  class ConstraintSet;
  class CounterCell;
  class DataRefObject;
  class Expr;
  class ExprSet;
  class Expression;
  class ExpressionSet;
  class FuncCallSite;
  class FuncCallSiteSet;
  class Interface;
  class InterfaceDefSet;
  class InterfaceVector;
  class InterfaceVectorSet;
  class Module;
  class ModuleDefSet;
  class ModulePort;
  class ModulePortSet;
  class NamedValue;
  class NamedValueSet;
  class NthExpr;
  class NthExprSet;
  class NthOperand;
  class NthOperandSet;
  class PackageDefSet;
  class PackageInstanceSet;
  class PackageInstanceVector;
  class PackageInstanceVectorSet;
  class PackageItem;
  class PackageItemSet;
  class PackageVector;
  class PackageVectorSet;
  class Program;
  class ProgramElement;
  class ProgramElementSet;
  class ProgramSet;
  class Scop;
  class ScopSet;
  class StringRefObject;
  class Structure;
  class StructureSet;
  class StructureItem;
  class StructureItemSet;
  class StructureInstance;
  class StructureInstanceSet;
  class StructureInstanceVector;
  class StructureInstanceVectorSet;
  class StructureMember;
  class StructureMemberSet;
  class StructureMemberVector;
  class StructureMemberVectorSet;
  class StructurePort;
  class StructurePortSet;
  class StructurePortVector;
  class StructurePortVectorSet;
  class Template;
  class TemplateSet;
  class TemplateValue;
  class TemplateValueSet;
  class TemplateVector;
  class TemplateVectorSet;
  class Type;
  class TypeSet;
  class Variable;
  class VariableSet;
  class VariableReference;
  class VariableReferenceSet;
  class Value;
  class ValueSet;
  class ValueVector;
  class ValueVectorSet;

  /*!
    \class VerilogPrinter
    \brief Printer for Verilog language.
  */
  class VerilogPrinter : public GenPrinter {
  public:
    /*!
      \brief Constructor.
    */
    VerilogPrinter();

    /*!
      \brief Destructor.
    */
    virtual ~VerilogPrinter();

    /*!
      \brief Start a new line.

      \return Value indicating success or failure.
    */
    bool StartNewLine();

    /*!
      \brief Finish a line.

      \return Value indicating success or failure.
    */
    bool FinishLine();

    /*!
      \brief Print a newline and indentation level.

      \return Value indicating success or failure.
    */
    bool PrintIndent();

    /*!
      \brief Print multiple newlines.

      \return Value indicating success or failure.
    */
    bool PrintNewLines(uint32_t aCount);

    /*!
      \brief Print a Verilog type.

      \return Value indicating success or failure.
    */
    bool PrintType(const Type* aType);

    /*!
      \brief Print a Verilog expression.

      \return Value indicating success or failure.
    */
    bool PrintExpr(const Expr* aExpr);

    /*!
      \brief Print a Verilog NthExpr.

      \return Value indicating success or failure.
    */
    bool PrintNthExpr(const NthExpr* aNthExpr);

    /*!
      \brief Print a Verilog Struct Instance.

      \param aInstance
      \param aStructure
      \