```verilog
module latch (input d, c, output wire [7:0] q, q_b );
wire [7:0] q_temp;