parameter NFIELDS = 32;
reg [0:NFIELDS-1] Result;