module test;
pack mypack;
reg mypack.x