```verilog
module tstdlatch