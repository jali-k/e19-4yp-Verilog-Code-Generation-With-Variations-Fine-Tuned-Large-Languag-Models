module Anding (input [1:0] a, b, output y);
endmodule
### Final Code: