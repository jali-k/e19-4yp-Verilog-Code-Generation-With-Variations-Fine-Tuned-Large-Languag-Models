module alu_mod(s, A, B, F);
input [2:0] s