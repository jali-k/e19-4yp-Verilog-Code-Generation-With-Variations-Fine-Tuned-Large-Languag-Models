module and2 (
input wire in_x,
input wire in_y,
output reg out_z
);
assign out_z = in_x & in_y;
endmodule
## 3. OR Gate
###