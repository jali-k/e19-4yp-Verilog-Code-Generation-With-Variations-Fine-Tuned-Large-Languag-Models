module sw2led2 (
input wire [7:0] sw,
output wire