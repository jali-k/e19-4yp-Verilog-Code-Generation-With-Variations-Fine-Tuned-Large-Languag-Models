module IR ( input [0:1] A [0:3], input [0:1] B [0:3], input load, clk,
output reg [0:1] add_out, output reg [0:1] mult_out );
// Simple