package mixed_sim_package;
const logic [31:0] ROM_CONSTANT = 'b11111111_11111111_111111