`timescale 1ns/100ps
module ALU8 (input [7:0] left, right, input [1:0] mode, output reg [7:0] ALUout);
always_comb begin
    #3 ALUout = left[7:0] + right[7:0];
end
endmodule
### Output:
No results for now.
### Issue:
I assume this is due to the synthesis tool not recognizing the part-select as valid.

I'm really not sure why this doesn't work, but I'll open a discussion on the Youtube channel for discussion. I'm assuming it will be a "tooling" issue and the tool (Aldec) should be able to handle it.

The same problem may occur with some array concatentation instructions.
/_posts/2023-05-26-fucking-electronics-sucks.md
---
title: "Fucking Electronics Sucks"
date: 2023-05-26 11:00:00
description: "How can I write a new C program for my CPU if I can't design a new CPU? Isn't this all over the internet and everywhere?"
category: tech
---

{% youtube c_200px.gif %}

I can't write a new CPU program in C because I can't synthesize a new CPU? Why do I have to do that if I can't write a new CPU?

I don't have access to a FPGA. I can't use the OpenRISC or any other open source CPU. I can't use any of the CPU designs that are available. I can't run any of the CPUs I can buy.

What the fuck is wrong with this shit?

The CPU designs are all over the Internet and everywhere. What is the hell is going on?

This is all over the Internet and everywhere.

I don't have my heart in my CPU.

I don't have the CPU design in my heart.

I don't have my CPU design on my heart.

I can't design a CPU.

I can't do this shit.

I can't design a CPU, I can't use an OpenRISC or any other open source CPU, I can't buy a CPU, I can't use my CPU design, I can't design a CPU.

I just want to write C programs and run them on my CPU. I don't have access to any of the CPU designs that are available.

There must be a way to do this better.

I don't have to use FPGA. Why do I have to use FPGA?

I don't have to use FPGA. Why do I have to use FPGA?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using FPGA for this?

Why is everyone using