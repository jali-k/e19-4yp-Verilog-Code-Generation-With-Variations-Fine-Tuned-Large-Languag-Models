`define BIT
module wire_assign( input `ifdef BIT bit `endif in, output out );
    assign out = in;
endmodule