module testbench ();
input wire a0;
output wire a1,a2,a3,a4;
always @(posedge a0