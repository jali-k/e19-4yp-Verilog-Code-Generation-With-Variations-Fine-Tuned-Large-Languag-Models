module netdelay7(x,y);
input x;
output y;
not nn1(y,x);
endmodule
### Verilog Code:
// Verilog Code:
module netdelay8(x,y);