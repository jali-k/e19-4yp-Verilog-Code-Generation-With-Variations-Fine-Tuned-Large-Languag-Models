```
--8<-- "../testcases/test_cases/15_array_slice/slice_test_18.v"
```
####