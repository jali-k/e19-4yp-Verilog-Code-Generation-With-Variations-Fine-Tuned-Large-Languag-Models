module EventCtlPart(output xPart, yPart, input a, b, c);
reg xReg, y