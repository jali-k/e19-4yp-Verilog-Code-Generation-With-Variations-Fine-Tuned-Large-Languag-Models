module testbench ();
generate struct { rand bit my_rand; } data;
process data;
endmodule