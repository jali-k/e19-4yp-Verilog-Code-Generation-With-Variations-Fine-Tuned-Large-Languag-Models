module wire_assign( input in, output reg out );
    assign out = in;
endmodule