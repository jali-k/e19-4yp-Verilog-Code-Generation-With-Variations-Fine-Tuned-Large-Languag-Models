module func8(x1, x2, x3, f