module Chap1Counter (Clk, Reset,