gates4_4 U1(
.x(sw),
.and4_(ld[3]),
.or4_(ld[2]),
.xor4_(ld[1]),
.and4_4_(ld[0]),
.priority(pri_ld)
);