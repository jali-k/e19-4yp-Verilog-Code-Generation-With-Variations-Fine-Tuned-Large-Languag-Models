module t_Clock_Prog ();
wire clock;
wire Resetn;

initial #100 $finish;
Clock_Prog M1 (clk, Resetn);
endmodule
1.2.6.2.5.2.5.2.4.2.5.2.5.2.4.3.5.2.5.2.5.2.4.4.2.5.2.5.2.4.3.5.2.5.2.4.3.4.5.2.5.2.4.3.5.2.5.2.4.4.3.5.2.5.2.4.3.5.2.5.2.4.4.4.5.2.5.2.4.3.5.2.5.2.4.4.4.4.5.2.5.2.4.3.5.2.5.2.4.4.4.4.4.5.2.5.2.4.3.5.2.5.2.4.4.4.4.4.4.5.2.5.2.4.3.5.2.5.2.4.4.4.4.4.4.4.5.2.5.2.4.3.5.2.5.2.4.4.4.4.4.4.4.4.5.2.5.