```
always @(w0 or w1 or w2 or w3 or S)
    case (S)
        {2'b00..2'b01}: