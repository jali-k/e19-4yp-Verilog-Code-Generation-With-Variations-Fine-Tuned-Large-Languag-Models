module Counter(input clk, input rst, output reg [