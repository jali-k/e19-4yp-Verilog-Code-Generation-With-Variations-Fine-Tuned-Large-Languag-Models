module Johnson_Counter (count, enable, clock, reset);
output [3: 0] count;
input enable;
input clock, reset;
reg [3: 0] count;
generate
for (genvar i = 0; i <= 4; i++) begin
always @ (posedge clock, posedge reset)
if (reset == 1) count <= 0;
else if (enable)
case (count)
4'b0000,
4'b0001,
4'b0011,
4'b0111,
4'b1111,
4'b1110,
4'b1100,
4'b1000: count <= {count[2: 0], 1'b1};
default: count <= 0;
endcase
end
endgenerate
endmodule

// 
### Verilog Code:
module Johnson_Counter (count, enable, clock, reset);
wire [3: 0] count;
reg enable;
reg clock, reset;
Johnson_Counter M0 (count, enable, clock, reset);
initial #500 $finish;
initial begin clock = 0; forever #5 clock = ~clock; end
initial fork
join
endmodule