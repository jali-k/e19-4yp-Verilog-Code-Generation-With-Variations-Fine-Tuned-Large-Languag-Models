module reg