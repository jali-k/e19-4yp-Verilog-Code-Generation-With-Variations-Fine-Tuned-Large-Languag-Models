module add32(a, b, cout, sum);
input [7:0] a, b;
output cout, [31:0] sum;
wire [4:0] a3;
wire [4:0] b3;
wire [4:0] a4;
wire [4:0] b4;
wire [4:0] a5;
wire [4:0] b5;
wire [4:0] a6;
wire [4:0] b6;
wire [4:0] a7;
wire [4:0] b7;
wire [4:0] a8;
wire [4:0] b8;
wire [4:0] a9;
wire [4:0] b9;
wire [4:0] a10;
wire [4:0] b10;
wire [4:0] a11;
wire [4:0] b11;
wire [4:0] a12;
wire [4:0] b12;
wire [4:0] a13;
wire [4:0] b13;
wire [4:0] a14;
wire [4:0] b14;
wire [4:0] a15;
wire [4:0] b15;
wire [4:0] a16;
wire [4:0] b16;
wire [4:0] a17;
wire [4:0] b17;
wire [4:0] a18;
wire [4:0] b18;
wire [4:0] a19;
wire [4:0] b19;
wire [4:0] a20;
wire [4:0] b20;
wire [4:0] a21;
wire [4:0] b21;
wire [4:0] a22;
wire [4:0] b22;
wire [4:0] a23;
wire [4:0] b23;
wire [4:0] a24;
wire [4:0] b24;
wire [4:0] a25;
wire [4:0] b25;
wire [4:0] a26;
wire [4:0] b26;
wire [4:0] a27;
wire [4:0] b27;
wire [4:0] a28;
wire [4:0] b28;
wire [4:0] a29;
wire [4:0] b29;
wire [4:0] a30;
wire [4:0] b30;
wire [4:0] a31;
wire [4:0] b31;
wire [4:0] a32;
wire [4:0] b32;
wire [4:0] a33;
wire [4:0] b33;
wire [4:0] a34;
wire [4:0] b34;
wire [4:0] a35;
wire [4:0] b35;
wire [4:0] a36;
wire [4:0] b36;
wire [4:0] a37;
wire [4:0] b37;
wire [4:0] a38;
wire [4:0] b38;
wire [4:0] a39;
wire [4:0] b39;
wire [4:0] a40;
wire [4:0] b40;
wire [4:0] a41;
wire [4:0] b41;
wire [4:0] a42;
wire [4:0] b42;
wire [4:0] a43;
wire [4:0] b43;
wire [4:0] a44;
wire [4:0] b44;
wire [4:0] a45;
wire [4:0] b45;
wire [4:0] a46;
wire [4:0] b46;
wire [4:0] a47;
wire [4:0] b47;
wire [4:0] a48;
wire [4:0] b48;
wire [4:0] a49;
wire [4:0] b49;
wire [4:0] a50;
wire [4:0] b50;
wire [4:0] a51;
wire [4:0] b51;
wire [4:0] a52;
wire [4:0] b52;
wire [4:0] a53;
wire [4:0] b53;
wire [4:0] a54;
wire [4:0] b54;
wire [4:0] a55;
wire [4:0] b55;
wire [4:0] a56;
wire [4:0] b56;
wire [4:0] a57;
wire [4:0] b57;
wire [4:0] a58;
wire [4:0] b58;
wire [4:0] a59;
wire [4:0] b59;
wire [4:0] a60;
wire [4:0] b60;
wire [4:0] a61;
wire [4:0] b61;
wire [4:0] a62;
wire [4:0] b62;
wire [4:0] a63;
wire [4:0] b63;
wire [4