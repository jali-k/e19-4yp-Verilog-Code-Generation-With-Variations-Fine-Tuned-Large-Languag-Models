module tst_nm_in();
  reg in; wire out;