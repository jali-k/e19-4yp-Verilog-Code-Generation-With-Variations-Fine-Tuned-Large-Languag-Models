module tb;
reg w0;
reg w1;
reg w2;
reg w3;
reg S;
reg f;