module test;
reg a, b, c;
assign b = 1;
assign c = 1;

always begin
    a = 1;
end

endmodule
##