module testbench ();
generate data;
  struct {
    rand bit [31:0] data;
  } data_struct;
process data;
endmodule