```
module mixed_sim;
reg dcontrol, x, y;
reg [31:0] data;
wire [31:0] bus;

package state_pkg;
reg [3:0] state_Mealy;
assign state_Mealy = {0,1,2,3,4,0,4,0};
always @(posedge state_Mealy[4])
begin
    case (state_Mealy[0])
        0:
            dcontrol = 1;
            data = 10;
        1:
            dcontrol = 1;
            data = 20;
        2:
            dcontrol = 1;
            data = 40;
        3:
            dcontrol = 0;
            data = 60;
    endcase
end
assign bus = dcontrol? data : 'bz;
always @(x)
y = ~x;
initial
begin
$monitor("time=%d dcontrol=%d data=%d x=%d y=%d bus=%d",
         $time, dcontrol, data, x, y, bus);
x = 1;
dcontrol = 0;
end
endmodule
```
### Result:
```
time=0 dcontrol=1 data=10 x=1 y=0 bus=10
time=1 dcontrol=1 data=20 x=0 y=1 bus=20
time=2 dcontrol=1 data=40 x=1 y=0 bus=40
time=3 dcontrol=0 data=60 x=0 y=1 bus=60
```
##### 2.2.2.2.3.2.2.3.2.4.2.5.2.6.2.7.2.8.1.2.3.3.2.2.2.3.2.2.3.3.2.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.1.2.3.3.2.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.2.2.3.3.1.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.3.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.4.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.5.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.6.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.7.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.8.2.3.9.2.2.3.10.2.2.3.11.9.2.3.10.2.2.3.11.10.2.3.11.2.2.3.11.11.2.3.11.3.2.3.11.4.2.3.11.5.2.3.11.6.2.3.11.7.2.3.11.8.2.3.11.9.2.3.11.10.1.2.3.3.2.3.4.2.3.5.2.3.6.2.3.7.2.3.8.2.3.9.2.3.10.2.3.11.2.3.11.3.2.3.11.4.2.3.11.5.2.3.11.6.2.3.11.7.2.3.11.8.2.3.11.9.2.3.11.10.2.3.11.11.
##### 2.2.2.2.3.2.2.3.4.1.2.3.5.2.2.3.6.1.2.3.7.1.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.1.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.1.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.1.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.2.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.3.2.3.4.2.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.4.2.3.5.2.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.5.2.3.6.2.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3.11.
##### 2.2.2.2.3.2.2.3.11.6.2.3.7.2.2.3.8.2.2.3.9.2.2.3.10.2.2.3