module tst_wand1;
reg i1,i2;
wire o;
wand1 ww(i1,i2,o);
always
begin
$display("i1=%b, i2=%b, o=%b",i1,i2,o);
if (((i1 >= 3'b0) && (i1 < 3'b1)) && ((i2 >= 3'b0) && (i2 < 3'b1))) begin o=3'b1; end
end
endmodule
### Expected Results:
i1=0, i2=0, o=0
i1=1, i2=0, o=0
i1=0, i2=1, o=0
i1=1, i2=1, o=1
### Observed Results:
i1=0, i2=0, o=0
i1=1, i2=0, o=0
i1=0, i2=1, o=0
i1=1, i2=1, o=1
```

## tst_wthres1

```
// Module: tst_wthres1
// Generated by LRM
// Description:
// Testbench for module wthres1.
//
// Note:
// 1. This testbench has 2 inputs, 1 output and 1 tristate.
// 2. The testbench generates 4 outputs, one for each input and three for
// the tristate.
// 3. The 4 outputs are compared to golden values to check for correctness.
//
// Usage:
// 1. Testbench parameters are read from the file tst_wthres1-params.txt.
// 2. The parameters file contains, one parameter per line.
// 3. The testbench can be started from the command prompt using the
// following syntax:
//  - "vcs -sverilog tst_wthres1.v -l vcs.log".
// 4. The simulator will generate a waveform of the testbench and its output.
// 5. Verilog/SystemVerilog code can be used to monitor the testbench.
// 6. After the test, the simulator will generate an output text file,
// "results.log", that contains all testbench outputs.
//
// Note: This testbench is not intended for synthesis.

`timescale 1ps / 1ps
// Testbench parameters are read from the file tst_wthres1-params.txt.
`include "tst_wthres1-params.txt"

// Source file: tst_wthres1.v
// Generated by LRM
// Description:
// Testbench for module wthres1.
//
// Note:
// 1. This testbench has 2 inputs, 1 output and 1 tristate.
// 2. The testbench generates 4 outputs, one for each input and three for
// the tristate.
// 3. The 4 outputs are compared to golden values to check for correctness.
//
// Usage:
// 1. Testbench parameters are read from the file tst_wthres1-params.txt.
// 2. The parameters file contains, one parameter per line.
// 3. The testbench can be started from the command prompt using the
// following syntax:
//  - "vcs -sverilog tst_wthres1.v -l vcs.log".
// 4. The simulator will generate a waveform of the testbench and its output.
// 5. Verilog/SystemVerilog code can be used to monitor the testbench.
// 6. After the test, the simulator will generate an output text file,
// "results.log", that contains all testbench outputs.
//
// Note: This testbench is not intended for synthesis.

`timescale 1ps / 1ps
// Testbench parameters are read from the file tst_wthres1-params.txt.
`include "tst_wthres1-params.txt"

// Source file: tst_wthres1.v
// Generated by LRM
// Description:
// Testbench for module wthres1.
//
// Note:
// 1. This testbench has 2 inputs, 1 output and 1 tristate.
// 2. The testbench generates 4 outputs, one for each input and three for
// the tristate.
// 3. The 4 outputs are compared to golden values to check for correctness.
//
// Usage:
// 1. Testbench parameters are read from the file tst_wthres1-params.txt.
// 2. The parameters file contains, one parameter per line.
// 3. The testbench can be started from the command prompt using the
// following syntax:
//  - "vcs -sverilog tst_wthres1.v -l vcs.log".
// 4. The simulator will generate a waveform of the testbench and its output.
// 5. Verilog/SystemVerilog code can be used to monitor the testbench.
// 6. After the test, the simulator will generate an output text file,
// "results.log", that contains all testbench outputs.
//
// Note: This testbench is not intended for synthesis.

`timescale 1ps / 1ps
// Testbench parameters are read from the file tst_wthres1-params.txt.
`include "tst_wthres1-params.txt"

// Source file: tst_wthres1.v
// Generated by LRM
// Description:
// Testbench for module wthres1.
//
// Note:
// 1. This testbench has 2 inputs, 1 output and 1 tristate.
// 2. The testbench generates 4 outputs, one for each input and three for
// the tristate.
// 3. The 4 outputs are compared to golden values to check for correctness.
//
// Usage:
// 1. Testbench parameters are read from the file tst_wthres1-params.txt.
// 2. The parameters file contains, one parameter per line.
// 3. The testbench can be started from the command prompt using the
// following syntax:
//  - "vcs -sverilog tst_wthres1.v -l vcs.log".
// 4. The simulator will generate a waveform of the testbench and its output.
// 5. Verilog/SystemVerilog code can be used to monitor the testbench.
// 6. After the test, the simulator will generate an output text file,
// "results.log", that contains all testbench outputs.
//
// Note: This testbench is not intended for synthesis.

`timescale 1ps / 1ps
// Testbench parameters are read from the file tst_wthres1-params.txt.
`include "tst_wthres1-params.txt"

// Source file: tst_wthres1.v
// Generated by LRM
// Description:
// Testbench for module wthres1.
//
// Note:
// 1. This testbench has 2 inputs, 1 output and 1 tristate.
// 2. The testbench generates 4 outputs, one for each input and three for
// the tristate.
// 3. The 4 outputs are compared to golden values to check for correctness.
//
// Usage:
// 1. Testbench parameters are read from the file tst_wthres1-params.txt.
// 2. The parameters file contains, one parameter per line.
// 3. The testbench can be started from the command prompt using the
// following syntax:
//  - "vcs -sverilog tst_wthres1.v -l vcs.log".
// 4. The simulator will generate a waveform of the testbench and its output.
// 5. Verilog/SystemVerilog code can be used to monitor the testbench.
// 6. After the test, the simulator will generate an output text file,
// "results.log", that contains all testbench outputs.
//
// Note: This testbench is not intended for synthesis.

`timescale 1ps / 1ps
// Testbench parameters are read from the file tst_wthres1-params.txt.
`include "tst_wthres1-params.txt"

// Source file: tst_wthres1.v
// Generated by LRM
// Description:
// Testbench for module wthres1.
//
// Note:
// 1. This testbench has 2 inputs, 1 output and 1 tristate.
// 2. The testbench generates 4 outputs