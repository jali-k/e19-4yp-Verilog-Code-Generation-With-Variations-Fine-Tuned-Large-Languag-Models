module Chap1Counter (Clk, Reset, Count);
input Clk,