# Generate a sequence of 1000 clock pulses
# Generate a reset pulse
# Generate a sequence of 1000 clock pulses

###