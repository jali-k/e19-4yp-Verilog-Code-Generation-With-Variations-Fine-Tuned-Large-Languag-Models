module netdelay6(x,y);
input x;
output y;
//assign y=x; // Assign 'x' to 'y' (direct assignment)
endmodule