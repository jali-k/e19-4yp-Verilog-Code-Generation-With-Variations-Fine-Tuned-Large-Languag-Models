module mux41b (
input wire [3:0] c,
input wire [1:0] s,
output wire z
);
assign z = ~s[1] & ~s[0] & c[0] // Select c[0] when s=00
| ~s[1] & s[0] & c[1] // Select c[1] when s=01
| s[1] & ~s[0] & c[2] // Select c[2] when s=10
| s[1] & s[0] & c[3]; // Select c[3] when s=11
| s[0] & s[1] & c[0] // Select c[0] when s=01
| s[0] & s[1] & c[1] // Select c[1] when s=10
| ~s[0] & ~s[1] & c[0] // Select c[0] when s=11
| ~s[0] & ~s[1] & c[1]; // Select c[1] when s=00
endmodule

### Code 1:

module mux81b(input wire [3:0] c,
input wire [1:0] s,
output wire z
);
wire [31:0] s1;
s1 = s;
s1[2] = s1[0];
assign z = ~s1[1] & ~s1[0] & c[0] // Select c[0] when s=00
| ~s1[1] & s1[0] & c[1] // Select c[1] when s=01
| s1[1] & ~s1[0] & c[2] // Select c[2] when s=10
| s1[1] & s1[0] & c[3]; // Select c[3] when s=11
| s1[0] & s1[1] & c[0] // Select c[0] when s=01
| s1[0] & s1[1] & c[1] // Select c[1] when s=10
| ~s1[0] & ~s1[1] & c[0] // Select c[0] when s=11
| ~s1[0] & ~s1[1] & c[1]; // Select c[1] when s=00
endmodule

### Code 2:

module mux81b(input wire [3:0] c,
input wire [1:0] s,
output wire z
);
wire [31:0] s1;
s1 = s;
s1[2] = s1[0];
assign z = ~s1[1] & ~s1[0] & c[0] // Select c[0] when s=00
| ~s1[1] & s1[0] & c[1] // Select c[1] when s=01
| s1[1] & ~s1[0] & c[2] // Select c[2] when s=10
| s1[1] & s1[0] & c[3]; // Select c[3] when s=11
| s1[0] & s1[1] & c[0] // Select c[0] when s=01
| s1[0] & s1[1] & c[1] // Select c[1] when s=10
| ~s1[0] & ~s1[1] & c[0] // Select c[0] when s=11
| ~s1[0] & ~s1[1] & c[1]; // Select c[1] when s=00

endmodule

### Input:

s=00, c=0000,0000,0000,0000,0000,0000,0000 // 0
s=00, c=0000,0000,0000,0000,0000,0000,0001 // 1
s=00, c=0000,0000,0000,0000,0000,0000,0010 // 2
s=00, c=0000,0000,0000,0000,0000,0000,0011 // 3
s=01, c=0000,0000,0000,0000,0000,0000,0000 // 4
s=01, c=0000,0000,0000,0000,0000,0000,0001 // 5
s=01, c=0000,0000,0000,0000,0000,0000,0010 // 6
s=01, c=0000,0000,0000,0000,0000,0000,0011 // 7
s=10, c=0000,0000,0000,0000,0000,0000,0000 // 8
s=10, c=0000,0000,0000,0000,0000,0000,0001 // 9
s=10, c=0000,0000,0000,0000,0000,0000,0010 // 10
s=10, c=0000,0000,0000,0000,0000,0000,0011 // 11
s=11, c=0000,0000,0000,0000,0000,0000,0000 // 12
s=11, c=0000,0000,0000,0000,0000,0000,0001 // 13
s=11, c=0000,0000,0000,0000,0000,0000,0010 // 14
s=11, c=0000,0000,0000,0000,0000,0000,0011 // 15

### Output:

s=00, c=0000,0000,0000,0000,0000,0000,0000 // 0
s=00, c=0000,0000,0000,0000,0000,0000,0001 // 1
s=00, c=0000,0000,0000,0000,0000,0000,0010 // 2
s=00, c=0000,0000,0000,0000,0000,0000,0011 // 3
s=01, c=0000,0000,0000,0000,0000,0000,0000 // 4
s=01, c=0000,0000,0000,0000,0000,0000,0001 // 5
s=01, c=0000,0000,0000,0000,0000,0000,0010 // 6
s=01, c=0000,0000,0000,0000,0000,0000,0011 // 7
s=10, c=0000,0000,0000,0000,0000,0000,0000 // 8
s=10, c=0000,00