```
inside
      {2{di}};
```
### Expected Output:
```
t=  20, clk=0, clr=0, pr=1, di=0, q=0 
t=  46, clk=0, clr=0, pr=0, di=0, q=0 
t=  48, clk=1, clr=1, pr=0, di=1, q=1 
t=  52, clk=0, clr=1, pr=0, di=1, q=1 
t=  54, clk=1, clr=1, pr=0, di=0, q=0 
t=  58, clk=0, clr=1, pr=0, di=0, q=0 
t=  60, clk=1, clr=1, pr=0, di=1, q=1 
t=  64, clk=0, clr=1, pr=0, di=1, q=1 
t=  66, clk=1, clr=1, pr=0, di=0, q=0 
t=  70, clk=0, clr=1, pr=0, di=0, q=0 
t=  72, clk=1, clr=1, pr=0, di=1, q=1 
t=  76, clk=0, clr=1, pr=0, di=1, q=1 
t=  78, clk=1, clr=1, pr=0, di=0, q=0 
t=  82, clk=0, clr=1, pr=0, di=0, q=0 
t=  84, clk=1, clr=1, pr=0, di=1, q=1 
t=  88, clk=0, clr=1, pr=0, di=1, q=1 
t=  90, clk=1, clr=1, pr=0, di=0, q