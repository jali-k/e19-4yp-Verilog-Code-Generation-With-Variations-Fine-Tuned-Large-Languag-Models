```c
#include <stdio