Always @(*)
begin: ALU
    Result <= ArgA [31:0] + ArgB [31:0];
end
### Expected Results:
Testcase: [31:0] (0)
Testcase: [31:0] (2**32)
Testcase: [31:0] (-2**32)
Testcase: [31:0] (2**32-1)
Testcase: [31:0] (-2**32+1)
Testcase: [31:0] (+1)
Testcase: [31:0] (-1)
Testcase: [31:0] (2**31-1)
Testcase: [31:0] (-2**31+1)
Testcase: [31:0] (2**31)
Testcase: [31:0] (-2**31)
Testcase: [31:0] (2**30-1)
Testcase: [31:0] (-2**30+1)
Testcase: [31:0] (2**30)
Testcase: [31:0] (-2**30)
Testcase: [31:0] (2**29-1)
Testcase: [31:0] (-2**29+1)
Testcase: [31:0] (2**29)
Testcase: [31:0] (-2**29)
Testcase: [31:0] (2**28-1)
Testcase: [31:0] (-2**28+1)
Testcase: [31:0] (2**28)
Testcase: [31:0] (-2**28)
Testcase: [31:0] (2**27-1)
Testcase: [31:0] (-2**27+1)
Testcase: [31:0] (2**27)
Testcase: [31:0] (-2**27)
Testcase: [31:0] (2**26-1)
Testcase: [31:0] (-2**26+1)
Testcase: [31:0] (2**26)
Testcase: [31:0] (-2**26)
Testcase: [31:0] (2**25-1)
Testcase: [31:0] (-2**25+1)
Testcase: [31:0] (2**25)
Testcase: [31:0] (-2**25)
Testcase: [31:0] (2**24-1)
Testcase: [31:0] (-2**24+1)
Testcase: [31:0] (2**24)
Testcase: [31:0] (-2**24)
Testcase: [31:0] (2**23-1)
Testcase: [31:0] (-2**23+1)
Testcase: [31:0] (2**23)
Testcase: [31:0] (-2**23)
Testcase: [31:0] (2**22-1)
Testcase: [31:0] (-2**22+1)
Testcase: [31:0] (2**22)
Testcase: [31:0] (-2**22)
Testcase: [31:0] (2**21-1)
Testcase: [31:0] (-2**21+1)
Testcase: [31:0] (2**21)
Testcase: [31:0] (-2**21)
Testcase: [31:0] (2**20-1)
Testcase: [31:0] (-2**20+1)
Testcase: [31:0] (2**20)
Testcase: [31:0] (-2**20)
Testcase: [31:0] (2**19-1)
Testcase: [31:0] (-2**19+1)
Testcase: [31:0] (2**19)
Testcase: [31:0] (-2**19)
Testcase: [31:0] (2**18-1)
Testcase: [31:0] (-2**18+1)
Testcase: [31:0] (2**18)
Testcase: [31:0] (-2**18)
Testcase: [31:0] (2**17-1)
Testcase: [31:0] (-2**17+1)
Testcase: [31:0] (2**17)
Testcase: [31:0] (-2**17)
### Actual Results:
Testcase: [31:0] (0)
Testcase: [31:0] (-2**32)
Testcase: [31:0] (2**32)
Testcase: [31:0] (-2**32+1)
Testcase: [31:0] (2**32-1)
Testcase: [31:0] (1)
Testcase: [31:0] (-1)
Testcase: [31:0] (-2**31+1)
Testcase: [31:0] (2**31-1)
Testcase: [31:0] (2**31)
Testcase: [31:0] (-2**31)
Testcase: [31:0] (-2**30+1)
Testcase: [31:0] (2**30-1)
Testcase: [31:0] (2**30)
Testcase: [31:0] (-2**30)
Testcase: [31:0] (-2**29+1)
Testcase: [31:0] (2**29-1)
Testcase: [31:0] (2**29)
Testcase: [31:0] (-2**29)
Testcase: [31:0] (-2**28+1)
Testcase: [31:0] (2**28-1)
Testcase: [31:0] (2**28)
Testcase: [31:0] (-2**28)
Testcase: [31:0] (-2**27+1)
Testcase: [31:0] (2**27-1)
Testcase: [31:0] (2**27)
Testcase: [31:0] (-2**27)
Testcase: [31:0] (-2**26+1)
Testcase: [31:0] (2**26-1)
Testcase: [31:0] (2**26)
Testcase: [31:0] (-2**26)
Testcase: [31:0] (-2**25+1)
Testcase: [31:0] (2**25-1)
Testcase: [31:0] (2**25)
Testcase: [31:0] (-2**25)
Testcase: [31:0] (-2**24+1)
Testcase: [31:0] (2**24-1)
Testcase: [31:0] (2**24)
Testcase: [31:0] (-2**24)
Testcase: [31:0] (-2**23+1)
Testcase: [31:0] (2**23-1)
Testcase: [31:0] (2**23)
Testcase: [31:0] (-2**23)
Testcase: [31:0] (-2**22+1)
Testcase: [31:0] (2**22-1)
Testcase: [31:0] (2**22)
Testcase: [31:0] (-2**22)
Testcase: [31:0] (-2**21+1)
Testcase: [31:0] (2**21-1)
Testcase: [31:0] (2**21)
Testcase: [31:0] (-2**21)
Testcase: [31:0] (-2**20+1)
Testcase: [31: