### Base Verilog Code:
module tstha_9();
   reg a,b; wire s,ca;
   ha_9 hh(s,ca,a,b); // Instantiate HA with rise/fall path delays
   initial begin a=0;b=0; end
   always begin #5 a=1;b=0; #5 a=0;b=1; #5 a=1;b=1; #5 a=0;b=0; end
   initial $monitor($time, " a = %b, b = %b,out carry = %b, outsum = %b ",a,b,ca,s);
   initial #30 $stop;
endmodule

module tstha_9();
  reg a,b; wire s,ca;
  ha_9 hh(.CLK(CLK),s,ca,a,b); // Instantiate HA with rise/fall path delays
  initial begin a=0;b=0; end
  always begin #5 a=1;b=0; #5 a=0;b=1; #5 a=1;b=1; #5 a=0;b=0; end
  initial $monitor($time, " a = %b, b = %b,out carry = %b, outsum = %b ",a,b,ca,s);
  initial #30 $stop;
endmodule

```

## Demonstrate Signal Routing