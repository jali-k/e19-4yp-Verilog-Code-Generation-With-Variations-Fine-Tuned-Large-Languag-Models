```verilog
module dff(D, Clock, Q);