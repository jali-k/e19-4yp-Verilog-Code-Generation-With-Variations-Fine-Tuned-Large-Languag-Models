module tst_nand1; //testbench
reg i1,i2;
wire o; // Added