module Anding (input a, b, output y);
and (y, a, b);
endmodule