module example3_2(enable, reset, data, led