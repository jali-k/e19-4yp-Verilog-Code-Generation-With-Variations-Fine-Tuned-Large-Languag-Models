module gade(a,a1,b,c,b1,c1);
input b,c,b1,c1;
output gade_intf a,a1;
// Instantiate OR gate with inertial delay 3
or #3 gg1(a1.c1,c1,b1);
// Instantiate AND gate with rise=2, fall=1 inertial delay
and #(2,1) gg2(a.c,c,b);
endmodule