```verilog
module t