[Download](https://github.com/tuhin18/ic/blob/master/tst_alu1.v)

### Outputs:
[![image](https://user-images.githubusercontent.com/41342513/126123579-71b714f3-5360-4863-8021-461dcfd2a82a.png)](https://github.com/tuhin18/ic/blob/master/tst_alu1.png)