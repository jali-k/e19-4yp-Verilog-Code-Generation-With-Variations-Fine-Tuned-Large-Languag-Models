module ALU (output logic signed [3:0] Result, input logic signed [3:0] ArgA, ArgB, input Clk);
endmodule
### Modified Simulation Output:
### Signed Arithmetic (signed inputs)
Result: 5'bd10
ArgA: 5'b00010
ArgB: 5'b00100
### Unsigned Arithmetic (unsigned inputs)
Result: 5'b10100
ArgA: 5'b00010
ArgB: 5'b00100