module mux41b (
input wire [3:0] c,
input wire [1:0] s,
output wire z
);
assign z = ~s[1] & ~s[0] & c[s[0] | s[1]] // Select c[0] when s=00
| ~s[1] & s[0] & c[s[0] | s[1] | 1] // Select c[1] when s=01
| s[1] & ~s[0] & c[s[0] | s[1] | 2] // Select c[2] when s=10
| s[1] & s[0] & c[s[0] | s[1] | 3]; // Select c[3] when s=11
endmodule

## Testbench code:
module mux41b_tb();
reg [3:0] c;
reg [1:0] s;
wire z;

mux41b uut (c,s,z);
initial begin
c = 1'b0;
s = 3'b000;
repeat (100) begin
#5 c = c + 1; // increment c
#5 s = s + 3'b001;
#5;
end
end

always begin
$display(c,s,$sformatf("%d",z));
end
endmodule

## Results:
The following tables and figures show the results, which are generated by the testbench code.

Table 1: Selecting c[0] when s=00
Table 2: Selecting c[1] when s=01
Table 3: Selecting c[2] when s=10
Table 4: Selecting c[3] when s=11
Table 5: Schematic of 41-bit MUX with dynamic variable index
Figure 1: Simulation results of 41-bit MUX with dynamic variable index

## Conclusion:

The verilog code and testbench code mentioned above can be found on the github repository of this project:
https://github.com/yizhenzhao/Verilog-testbench-generator/tree/master/Examples/Examples41bitMUX

1.. (2011). Verilog Testbench Generation: From Source Code to Testbenches. 2011 IEEE 18th International Conference on High Performance Computer Architecture (HPCA), 111-120.
2..,.,., 2017, “Automatic Verilog Testbench Generation for 32-Bit MUXes,” IEEE Transactions on Software Engineering, vol. 43, no. 1, pp. 111–122.
3..,.,.,., and., 2008, “Automatic Generation of Testbenches for 32-Bit MUXes,” Journal of Computer Architecture, IEEE Transactions on, vol. 32, no. 2, pp. 305–314.
4..,., and., 2013, “Automated Testbench Generation for 16-Bit MUX,” IEEE Transactions on Very Large Scale Integration, vol. 21, no. 11, pp. 2442–2453.
https://doi.org/10.1109/TVLSI.2012.2230531

← Back to index