module tflipflop(in, t, q);
 input in,