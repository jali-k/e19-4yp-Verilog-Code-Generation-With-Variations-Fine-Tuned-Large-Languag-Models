module full_adder_chain(B, B_R, Cin, S, Cout);
input B, B_R, Cin;
output S, Cout;

module full_adder_chain(B, B_R, Cin, S, Cout);

input B, B_R, Cin;
output S, Cout;

## 4.8 Designing the 4-Bit Binary Decoder

### Explanation:
4-Bit Binary Decoder is designed to input four bits and output four bits. It is an M-type gate with an invert gate. It is used