#include <stdio.h>
  #include <stdint.h>
  typedef struct { unsigned a; int b; } ha_1_t1;
  typedef struct