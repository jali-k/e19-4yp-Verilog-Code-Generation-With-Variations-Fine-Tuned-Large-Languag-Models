module EventCtlPart (output xPart, yPart, input a, b, c);
reg xReg, yReg;
assign xPart = xReg;
assign yPart = yReg;
always @(*)
begin: PartList
    xReg <= a & b & c;
    yReg <= (b | c) ^ a;
end
EventCtlPart #(.Range(2),.Slice(3)) 
endmodule
### Testbench Code:
module testbench;
reg a, b, c;
EventCtlPart e(a, b, c);
initial $dumpfile("x.vcd");
initial
$dumpvars(0, e);
initial #10;
a <= 1;
b <= 1;
c <= 0;
initial #10;
a <= 1;
b <= 1;
c <= 1;
initial #10;
a <= 1;
b <= 0;
c <= 1;
initial #10;
a <= 0;
b <= 1;
c <= 1;
initial #10;
a <= 0;
b <= 0;
c <= 1;
initial #10;
a <= 0;
b <= 0;
c <= 0;
initial #10;
a <= 1;
b <= 0;
c <= 0;
initial #10;
a <= 1;
b <= 1;
c <= 0;
initial #10;
a <= 0;
b <= 1;
c <= 0;
initial #10;
a <= 0;
b <= 0;
c <= 0;
#10;
$finish;
endmodule
# Copyright (c) 2013-2014,  ()
# Released under the 2-clause BSD license (see the file LICENSE for details)

all: test

test: run_test.py test_data
	python run_test.py

test_data: test_data.py
	python test_data.py

clean:
	rm -rf *.pyc __pycache__
.. _section-1:

Getting started
===============

After installing VUnit, you can start writing your first test.

It is recommended to write your own tests following the `PEP8 <http://www.python.org/dev/peps/pep-0008/>`_ rules. This will make your code easier to read and maintain.

Here is a simple example which creates two test modules, ``test_module1`` and ``test_module2``, each containing one test:

.. code-block:: python

    from vunit import VUnit
    from vunit.utils import Test

    VUnit.add_class_path(r"C:\MySource\my_unit")
    VUnit.add_class_path(r"C:\MySource\my_unit2")

    @VUnit.main()
    def main():
        # Create instances of the modules to be tested
        module1 = Test(r"my_unit.test_module1")
        module2 = Test(r"my_unit2.test_module2")
   
        # Create the testbench with the modules to be tested
        tb = Test.create(module1)
        Test.create(module2)

        # Run the testbench
        tb.run()

    if __name__ == "__main__":
        main()

If you save the above script as ``my_test.py``, you can now run it with the command:

.. code-block:: bash

    $ python my_test.py

This should create a new directory named ``__vunit_output__`` in the same directory that ``my_test.py`` resides in, containing the following files:

* ``my_test.out``: The output of the simulation with VUnit
* ``my_test.log``: The log file created by VUnit
* ``my_test.vcd``: The VCD file generated by the simulation

This is what ``my_test.out`` contains:

.. code-block:: text

    +--------------------------------------------------------------+
    | Summary                                                     |
    +--------------------------------------------------------------+
    | test_module1.test_case_1                                    |
    |                                                               |
    | Finished in 0.000 s                                          |
    |                                                               |
    | Failures: 0                                                  |
    | Errors: 1                                                    |
    |                                                               |
    | Exit code: 0                                                 |
    |                                                               |
    +--------------------------------------------------------------+

It is possible to get more information about the failed test with the following command:

.. code-block:: bash

    $ python -m vunit.run_test -u -v my_test.py

This will create a new directory named ``__vunit_output__`` in the same directory that ``my_test.py`` resides in, containing the following files:

* ``my_test.out``: The output of the simulation with VUnit
* ``my_test.log``: The log file created by VUnit
* ``my_test.vcd``: The VCD file generated by the simulation
* ``my_test.summary``: The "detailed" report of the simulation
* ``my_test.errors``: The list of errors encountered during simulation

This is what ``my_test.errors`` contains:

.. code-block:: text

    +--------------------------------------------------------+-----------------+
    | Failure                                               |                 |
    +--------------------------------------------------------+-----------------+
    | my_unit.test_module1.test_case_1 > tb.module1.test    | My error message |
    +--------------------------------------------------------+-----------------+

You now know how to write your first tests!

.. toctree::
   :glob:
   :maxdepth: 1

   getting_started/examples/*
.. _section-1:

Getting started
===============

After installing VUnit, you can start writing your first test.

It is recommended to write your own tests following the `PEP8 <http://www.python.org/dev/peps/pep-0008/>`_ rules. This will make your code easier to read and maintain.

Here is a simple example which creates two test modules, ``test_module1`` and ``test_module2``, each containing the same test:

.. code-block:: python

    from vunit import VUnit
    from vunit.utils import Test

    VUnit.add_class_path(r"C:\MySource\my_unit")
    VUnit.add_class_path(r"C:\MySource\my_unit2")

    @VUnit.main()
    def main():
        # Create instances of the modules to be tested
        module1 = Test(r"my_unit.test_module1")
        module2 = Test(r"my_unit2.test_module2")
   
        # Create the testbench with the modules to be tested
        tb = Test.create(module1)
        Test.create(module2)

        # Run the testbench
        tb.run()

    if __name__ == "__main__":
        main()


You now know how to write your first tests!

.. toctree::
   :glob:
   :maxdepth: 1

   getting_started/examples/*
import pytest
from vunit import VUnit


@pytest.fixture(scope="session", autouse=True)
def setup_vunit():
    VUnit.add_class_path(".")
    VUnit.add_class_path("../../../test_data/test_module")
    VUnit.add_class_path("../../../test_data/test_module/mod")
    VUnit.add_class_path("../../../test_data/test_module/mod2")
    VUnit.add_class_path("../../../test_data/sub_module")
    VUnit.add_class_path("../../../test_data/sub_module/mod3")
# Copyright (c) 2013-2014,  ()
# Released under the 2-clause BSD license (see the file LICENSE for details)

import os
import sys
from shutil import rmtree
from zipfile import ZipFile

from vunit.test_suite import Test
from vunit.cli import run_cli

try:
    import pytest
except ImportError:
    def pytest_collect_file(parent, path):
        return None

try:
    from StringIO import StringIO
except:
    from io import StringIO


def pytest_addoption(parser):
    parser.addoption(
        "--test_folder",
        action="store",
        help="Specify the folder to be used as test folder",
    )
    parser.addoption(
        "--test_module",
        action="store",
        help="Specify the name of the test module",
    )


def pytest_report_header(config):
    if config.getoption("--test_module"):
        return "Run test: {} {}".format(config.getoption("--test_module"),
                                        config.getoption("--test_folder"))


def pytest_cmdline_main(config):
    run_cli()