module Prob_6_7_Mealy (Detect_Mealy, di, clk, rst);
// Mealy nonresetting sequence detector
output Detect_Mealy;
input di, clk, rst;
parameter S_0 = 0, S_1 = 1, S_2 = 2, S_3 = 3;
parameter S_5 = 5, S_6 = 6, S_7 = 7;
reg [2: 0] state_Mealy, next_state;
wire Detect_Mealy = (((state_Mealy == S_3)&&(di$inside$0))|((state_Mealy == S_7)&&(di$inside$1))); always @ (posedge clk) if (rst) state_Mealy <= S_0; else state_Mealy <= next_state; always @ (state_Mealy, di) begin next_state = S_0; case (state_Mealy) S_0: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_5; S_1: if (di$inside$0) next_state = S_2; else if (di$inside$1) next_state = S_5; S_2: if (di$inside$0) next_state = S_3; else if (di$inside$1) next_state = S_5; S_3: if (di$inside$0) next_state = S_3; else if (di$inside$1) next_state = S_5; S_5: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_6; S_6: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_7; S_7: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_7; default: next_state = S_0; endcase end always @ (posedge clk) if (rst) state_Mealy <= S_0; else state_Mealy <= next_state; endmodule ### Variation Instruction: In the behavioral D-latch, use `inside` operator on `di` to check against a single-bit value of a fixed array slice. ### Modified Code: module Prob_6_7_Mealy (Detect_Mealy, di, clk, rst); // Mealy nonresetting sequence detector output Detect_Mealy; input di, clk, rst; parameter S_0 = 0, S_1 = 1, S_2 = 2, S_3 = 3; parameter S_5 = 5, S_6 = 6, S_7 = 7; reg [2: 0] state_Mealy, next_state; wire Detect_Mealy = (((state_Mealy == S_3)&&(di$inside$0))|((state_Mealy == S_7)&&(di$inside$1))); always @ (posedge clk) if (rst) state_Mealy <= S_0; else state_Mealy <= next_state; always @ (state_Mealy, di) begin next_state = S_0; case (state_Mealy) S_0: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_5; S_1: if (di$inside$0) next_state = S_2; else if (di$inside$1) next_state = S_5; S_2: if (di$inside$0) next_state = S_3; else if (di$inside$1) next_state = S_5; S_3: if (di$inside$0) next_state = S_3; else if (di$inside$1) next_state = S_5; S_5: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_6; S_6: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_7; S_7: if (di$inside$0) next_state = S_1; else if (di$inside$1) next_state = S_7; default: next_state = S_0; endcase end always @ (posedge clk) if (rst) state_Mealy <= S_0; else state_Mealy <= next_state; endmodule ## Problem 7: Mealy NonResetting Moore Sequence Detector ### Base Verilog Code: module Prob_7_moore_nr (Detect_moore_nr, D_in, clk, rst); // Nonresetting moore sequence detector output Detect_moore_nr; parameter S_0 = 0, S_1 = 1, S_2 = 2, S_3 = 3; parameter S_10 = 10, S_11 = 11, S_12 = 12, S_13 = 13; input D_in, clk, rst; reg [2: 0] state_moore_nr, next_state; wire Detect_moore_nr = (((state_moore_nr == S_3)&&(D_in == 0))|((state_moore_nr == S_13)&&(D_in == 1))); always @ (posedge clk) if (rst) state_moore_nr <= S_0; else state_moore_nr <= next_state; always @ (D_in, clk) begin next_state = S_0; case (D_in) S_0: next_state = S_1; S_1: next_state = S_2; S_2: if (state_moore_nr == S_3) next_state = S_3; else if (state_moore_nr == S_13) next_state = S_13; S_3: if (state_moore_nr == S_3) next_state = S_3; else if (state_moore_nr == S_13) next_state = S_13; S_13: if (state_moore_nr == S_3) next_state = S_3; else if (state_moore_nr == S_13) next_state = S_13; default: next_state = S_0; endcase end always @ (posedge clk) if (rst) state_moore_nr <= S_0; else state_moore_nr <= next_state; endmodule ### Variation Instruction: In the behavioral D-latch, use `inside` operator on `di` to check against a fixed array slice from a dollar unit constant. ### Modified Code: module Prob_7_moore_nr (Detect_moore_nr, di, clk, rst); // Nonresetting moore sequence detector output Detect_moore_nr; input di, clk, rst; parameter S_0 = 0, S_1 = 1, S_2 = 2, S_3 = 3; parameter S_10 = 10, S_11 = 11, S_12 = 12, S_13 = 13; reg [2: 0] state_moore_nr, next_state; wire Detect_moore_nr = (((state_moore_nr == S_3)&&(di$inside$0))|((state_moore_nr == S_13)&&(di$inside$1))); always @ (posedge clk) if (rst) state_moore_nr <= S_0; else state_moore_nr <= next_state; always @ (D_in, clk) begin next_state = S_0; case (D_in) S_0: next_state = S_1; S_1: next_state = S_2; S_2: if (state_moore_nr == S_3) next_state = S_3; else if (state_moore_nr == S_13) next_state = S_13; S_3: if (state_moore_nr == S_3) next_state = S_3; else if (state_moore_nr == S_13) next_state = S_13; S_13: if (state_moore_nr == S_3) next_state = S_3; else if (state_moore_nr == S_13) next_state = S_13; default: next_state = S_0; endcase end always @ (