module clock_gen_forever;
  reg clk;
  initial clk=1'b0;
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("clk=%b, t=%0d", clk,$time);
  initial #2 $monitor("