### Variation Description:
Add a parameter called N to the module declaration. The parameter specifies how large the output port should be. In the module body, generate the output port as a N-bit output port.
### Variation Inst