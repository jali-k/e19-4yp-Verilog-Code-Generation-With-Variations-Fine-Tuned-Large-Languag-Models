```Verilog
module program(F, R);
input [3:0] F;
output reg [3:0] R;

endmodule
```
### Explanation:
`F[3:0]` are the `inputs` of the module. The `R` is the result of the module.

## Testbenches
The testbench for the `program` module will be a normal testbench with 8 testcases.

### Testcase1:
The testcase1 will be a test with all values of `F`.

### Testcase2:
The testcase2 will be a test with all values of `F`.

### Testcase3:
The testcase3 will be a test with all values of `F`.

### Testcase4:
The testcase4 will be a test with all values of `F`.

### Testcase5:
The testcase5 will be a test with all values of `F`.

### Testcase6:
The testcase6 will be a test with all values of `F`.

### Testcase7:
The testcase7 will be a test with all values of `F`.

### Testcase8:
The testcase8 will be a test with all values of `F`.

# The `program_tb` testbench

The `program_tb` testbench is a testbench that will test the functionality of the `program` module. It will be a normal testbench with 8 testcases. The testcases will be the following:

### Testcase1: 
The testcase1 will be a test with all values of `F`.

### Testcase2:
The testcase2 will be a test with all values of `F`.

### Testcase3:
The testcase3 will be a test with all values of `F`.

### Testcase4:
The testcase4 will be a test with all values of `F`.

### Testcase5:
The testcase5 will be a test with all values of `F`.

### Testcase6:
The testcase6 will be a test with all values of `F`.

### Testcase7:
The testcase7 will be a test with all values of `F`.

### Testcase8:
The testcase8 will be a test with all values of `F`.

# The `main_tb` testbench

The `main_tb` testbench is a testbench that will test the functionality of the modules that will be used to build the chip. It will be a normal testbench with 8 testcases. The testcases will be the following:

### Testcase1: 
The test