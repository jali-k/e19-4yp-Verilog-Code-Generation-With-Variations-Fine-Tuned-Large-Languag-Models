```
struct randval {
 int rand;
};

module testbench ();
generate data;
process data;
endmodule
### Output:

```
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 6
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 0 ns
Description: 
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 0 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 0 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 0 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 15168
Thread ID (TID): 15168
File: /home/yousef/Desktop/Veri-Random/src/testbench.v
Line: 7
Name: TESTBENCH_TOP
Module: testbench
Clock: 500000
State: Running
Time: 1 ns
Description: Generate statement: for (i=0; i<10; i=i+1)
== Testbench ==
Process ID (PID): 151