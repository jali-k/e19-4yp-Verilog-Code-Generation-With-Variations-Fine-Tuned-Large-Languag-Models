```verilog
module mealy