```

```verilog
### Base Verilog Code: