initial
    in =1'b1; // Start with input high -> output low
  always
  initial $monitor($time, " in = %b, output = %b ",in,out);
  initial #15 $stop; // Stop simulation
endmodule
### Result:
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1, output =  0
in =  1