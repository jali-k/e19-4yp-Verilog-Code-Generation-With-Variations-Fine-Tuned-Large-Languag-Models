```
index = inside(index, 0, 1, 2, 3, 4, 5, 6, 7);
```
### Previous Counter Instantiation:
```
jk ff[7:0](clk, reset, j, k, q, qbar, index[0], index[1], index[2], index[3], index[4], index[5], index[6], index[7]);
```
### Modified Counter Instantiation:
```
jk ff[7:0](clk, reset, j, k, q, qbar, index[0], index[1], index[2], index[3], index[4], index[5], index[6], index[7]);
```
### Counter Outputs:
<img width="234" alt="Screen Shot 2023-03-07 at 9 51 10 PM" src="https://user-images.githubusercontent.com/66631285/223611469-d59a73e0-97e0-4e91-aa7d-7320d28d55b7.png">


### Logic Diagram:
![Screen Shot 2023-03-07 at 9 51 38 PM](https://user-images.githubusercontent.com/66631285/223611664-11322e94-904f-485e-812c-6bba59cbf483.png)