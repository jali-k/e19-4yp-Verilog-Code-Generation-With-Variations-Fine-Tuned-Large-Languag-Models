module aoibeh2(o,a,b); // Mixed structural/behavioral AOI
output o;
input[1:0]a,b;
wire a1,b1; // Outputs of AND gates
wire f1; // Outputs of OR gate
reg o; // Behavioral output must