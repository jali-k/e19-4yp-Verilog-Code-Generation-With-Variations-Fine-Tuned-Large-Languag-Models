assign Output = InputA*InputB;

### Changes:

1) The wire type Output has been changed to