```
initial begin: Apply_Data
generate
for (indx=0; indx<8