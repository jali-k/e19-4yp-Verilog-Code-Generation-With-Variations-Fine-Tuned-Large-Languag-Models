1) module ALU ( input [7:0] a, b, input pass, add,
2) output logic[7:0] alu_out );