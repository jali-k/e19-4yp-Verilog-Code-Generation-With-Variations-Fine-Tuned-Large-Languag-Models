
module top
(
  input CLK,
  input RST,
  output [7:0] led
);

  assign led = 8;

endmodule
