module tb_TOP1;
  reg CLK, RST_X;
  wire [1:0] x_comparator;
  wire [1:0] y_comparator;
  wire [1:0] z_comparator;
  wire [1:0] p_comparator;
  wire [1:0] q_comparator;
  wire [1:0] r_comparator;
  wire [1:0] s_comparator;
  wire [1:0] t_comparator;
  wire [1:0] u_comparator;
  wire [1:0] v_comparator;
  wire [1:0] w_comparator;
  wire [1:0] x_comparator;
  wire [1:0] y_comparator;
  wire [1:0] z_comparator;
  TOP1 uut(.CLK(CLK),.RST_X