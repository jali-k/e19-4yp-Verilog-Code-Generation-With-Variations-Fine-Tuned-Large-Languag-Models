module contres(o,i1,i2);
input i1,i2;
output o;
// Drive wire 'o' from two buffers with specified output strengths
buf(pull1, weak0) g1(o,i1); // Drives pull '1', weak '0'
buf(pull1, weak0) g2(o,i2); // Drives pull '1', weak '0'
// Resolution: 1,1->1; 1,0->1; 0,1->1; 0,0->0; 1,Z->1; 0,Z->X; Z,Z->Z
// Effective behavior is OR due to pull1 dominance over weak0
// Assign array values
assign i1 = {1'b0, 2'b10, 3'b0};
assign i2 = {i1[0], 1'b0};
assign o = i1[0] | i2[0];
i1 <= {1'b0, 2'b10, 3'b0}; // assign array values with <= operator
endmodule

## [4-23] Array Assignment with Assignment Operator (Alternate)

### Original Code:
module contres(o,i1,i2);
input i1,i2;
output o;
// Drive wire 'o' from two buffers with specified output