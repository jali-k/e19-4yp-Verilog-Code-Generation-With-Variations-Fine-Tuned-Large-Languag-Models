module dff(do,di,clk); // Behavioral D Flip-Flop
output do;
input di,clk;
reg do; // Output must be reg for procedural assignment
initial
do=1'b0; // Initialize output
// Assign input 'di' to output 'do' on negative clock edge
always@(negedge clk) do = di; // Use non-blocking <= for sequential logic
endmodule
The case statement can also be implemented in C style, i.e., without the need for the 'case' keyword.
### Base Verilog Code: