### Test Code:
### Verilog Code: