```verilog
module clock_gen_forever_with_function;
  reg clk, en;
  reg [3:0] counter;
  
  // Function to generate a random number
  function [3:0] generateRandomNumber;
    input [3:0] lastNumber;
    begin
      generateRandomNumber = lastNumber + ($random % 7); // Calculate a random number in range [lastNumber, lastNumber + 6]
    end
  endfunction
  
  // Generate clock using for loop, controlled by 'en'
  always @(posedge en) // Start clock generation on posedge en
    begin
      counter = generateRandomNumber(counter); // Use function to get a random counter value
      for (int i=0; i<counter; i++) // The number of times the loop runs is determined by the counter
      begin
        #2 clk = ~clk; // Toggle clock every 2 time units
      end
    end
  
  initial
  begin
    clk = 1'b0; // Initialize clock
    en = 1'b0; // Start disabled
    counter = 0; // Initialize counter to 0
  end
  
  initial $monitor("clk=%b, t=%0d, en=%b, counter=%0d", clk, $time, en, counter);
endmodule
```
This code will generate a clock with a random period between 2 to 8 time units. The random number generated by the function is stored in the `counter` register, and this value is used as the number of times the loop runs in the forever loop. The random number generated is in range [lastNumber, lastNumber + 6] inclusive. Each run of the loop will generate a new random number for the next run. 

Remember to put the `$monitor` back to the code if you intend to use this code for testing in a simulator. It is mainly used for debugging purposes.###

Note: The function `$random()` is used to generate a random number. The random number is between 0 and 32767 (2^15-1). The input and output of the function is of type `reg [3:0]`, which means