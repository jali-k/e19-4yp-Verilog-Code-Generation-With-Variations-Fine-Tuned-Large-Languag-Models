module latch (input d, c, output q, q_b );
always begin
wait ( c );
end
endmodule
1.
The behavior of the test-bench is the same as the Base Verilog.
2.
The Verilog-Source code is not synthesizable.
3.
The Verilog-Source code is synthesizable. However, the synthesized netlist cannot be implemented in either Xilinx or Altera.
4.
The Verilog-Source code is synthesizable. The synthesized netlist can be implemented in both Xilinx and Altera.
5.
None of the above.

## 5.
A test-bench is required to test a Verilog-Source code, but only test-benches are not sufficient. A test-bench must also include a test-vector.
1.
True
2.
False
3.
None of the above

## 6.
A test-bench must include a test-vector in order to test a Verilog-Source code.
1.
True
2.
False
3.
None of the above

## 7.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
0
0
1
0
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
0
0
1
0
1
1
1
0
0
1
0
1
0
1
0
1
0
1
1
1
1
1
1
1
1
1

## 8.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 9.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 10.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 11.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 12.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 13.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 14.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 15.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 16.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 17.
The test-vector for the latch is the following:
d
c
q
q_b
1
1
1
1
0
1
1
0
1
0
1
1
1
0
1
1
1
1
0
1
1
0
1
1
1
0
1
1
0
1
1
1
1
1
1
1
1
1

## 18.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 19.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 20.
The test-vector for the latch is the following:
d
c
q
q_b
0
0
0
0
1
0
0
1
1
1
1
0
0
1
1
1
0
0
1
0
1
1
1
0
1
1
0
1
0
1
1
1
1
1
1
1
1
1

## 21.
The test-vector for the latch is the following:
d
c
q
q_b
1
1
1
1
0
1
1
0
1
0
1
1
1
0
1
1
1
1
0
1
1
0
1
1
1
0
1
1
0
1
1
1
1
1
1
1
1
1

## 22.
The test-vector for the latch is the following:
d
c
q
q_b
1
1
1
1
0
1
1
0
1
0
1
1
1
0
1
1
1
1
0
1
1
0
1
1
1
0
1
1
0
1
1
1
1
1
1
1
1
1

## 23.
The test-vector for the latch is the following:
d
c
q
q_b
1
1
1
1
0
1
1
0
1
0
1
1
1
0
1
1
1
1
0
1
1
0
1
1