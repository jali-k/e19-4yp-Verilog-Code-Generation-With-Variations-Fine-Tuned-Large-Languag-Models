module EventCtlPart_v2 (output xPart, yPart, input a, b, c);

reg xReg, yReg;
assign xPart = xReg;
assign yPart = yReg;

always @(a,b)
begin: PartList
    xReg <= a & b & c;
    yReg <= (b | c) ^ a;
end
endmodule

### Generated Verilog:
module EventCtlPart_v2 (output xPart, yPart, input a, b, c);
    reg xReg, yReg;
    output xPart;
    output yPart;
    input a;
    input b;
    input c;
    always @(a,b) begin: PartList
        xReg <= a & b & c;
        yReg <= (b | c) ^ a;
    end
endmodule

### Results:
The original code has a more straightforward flow, but the Verilog generated by it is longer as it requires a 2D to represent all 8 nested ifs. The modified version uses a 3D array to represent the 8 different branching possibilities. This is not as clear on the flow, but simplifies the Verilog code.
### Notes:
I am not sure if the modified code is correct. I tried to simplify it to an array of 32 elements. The array index was determined using a 2 bit variable. But I couldn't use a 3 bit variable. The 3 bit variable is not supported in System Verilog.
#include "EventCtlPart_v2.h"
#include <iostream>

//int main()
int main(int argc, char* argv[])
{
    std::vector<EventCtlPart_v2*> instances;
    char ch;
    int a, b, c;
    do {
        std::cout << "Enter a, b, c values:";
        std::cin >> a >> b >> c;
        std::cout << "Create a new instance? (y/n):";
        std::cin >> ch;
        
        EventCtlPart_v2* part;
        
        if ((ch == 'y') || (ch == 'Y'))
        {
            part = new EventCtlPart_v2;
            instances.push_back(part);
        }
       ut << part->xPart << " | " << part->yPart << std::endl;
        }   
    } while (ch == 'y' || ch == 'Y');
}
 
        if (part!= NULL)
        {
            part->a = a;
            part->b = b;
            part->c = c;
            
            std::co:
	g++ -c EventCtlPart.cpp

EventCtlPart_v2.o: EventCtlPart_v2.cpp EventCtlPart_v2.h
	g++ -c EventCtlPart_v2.cpp

main.o: main.cpp
	g++ -c main.cpp

clean:
	rm *.o
EventCtlPart: EventCtlPart.o EventCtlPart_v2.o main.o
	g++ -o EventCtlPart EventCtlPart.o EventCtlPart_v2.o main.o

EventCtlPart.o