module Prob_9 (Detect, D_in, clk, rst);
// D flipflop with edge detector
output Detect;
input D_in, clk, rst;