module t_John