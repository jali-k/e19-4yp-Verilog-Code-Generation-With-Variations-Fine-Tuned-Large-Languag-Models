```
logic [7:0] a;               // variable declaration
logic [7:0] b;
logic [7:0] c;
  initial begin
        a = {8{1'b0}};  // initialization of a
        b = {8{1'b0}};  // initialization of b
        c = {8{1'b1}};  // initialization of c
    end
```

### Differences


### Conclusion:



### References:
[1] [Verilog Initialization](https://verilog.as/2018/10/11/verilog-initializations.html)
[2] [Verilog Initialization](https://www.doulos.com/knowhow/verilog/initialization/)
[3] [Verilog Initialization](https://github.com/HandsOnOpenSource/Verilog-Coding-Standard/blob/master/Verilog%20Initialization.md)