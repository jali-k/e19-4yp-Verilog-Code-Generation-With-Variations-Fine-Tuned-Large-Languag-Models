module gbe(a,b,c,d,e,f,