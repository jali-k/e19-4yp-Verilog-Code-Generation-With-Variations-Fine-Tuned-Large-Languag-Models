module CMOSsw1(output reg