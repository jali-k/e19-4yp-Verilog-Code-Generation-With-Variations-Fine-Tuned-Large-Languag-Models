module ttst_ttrimux2_1(); // Assuming this tests a tristate 2-to-1 mux called ttrimux2_1
reg e;
reg [1:0]i; // Should be reg i0, i1; or reg [0:0] i0, i1; or just input wires if MUX takes separate inputs
reg s;
wire out; // Added wire declaration
// ttrimux2_1 mm(out,e,i,s); // Instantiation requires correct MUX definition
initial
begin
e =0; i = 2'b00; s = 1'b0; // Added initial's' value
end
always
begin
end
generate
begin
initial $monitor($time," enable e = %b, s= %b, input i = %b,output out = %b ",e,s,i,out); end endmodule ### Result ### Before: enable e = 0, s= 0, input i = 00,output out = 0 In the original testbench, the enable was being set to 0 in the initial block before the test began. This caused the same result in the sliced output as it did in the DUT. ### After: enable e = 0, s= 0, input i = 00,output out = 0 In the modified testbench, the enable was being set to 0 in the initial block before the test began. This caused the same result in the sliced output as it did in the DUT. However, after the enable was replaced with the generate block, the enable was set to 1 in the initial block because the generate block sets s to 1'b1. This caused a different result in the sliced output. ### Conclusion: The reason the enable was not being reset to 0 in the generate block was because it was not being set using a generate statement. In the original testbench, it was being set using a statement in the initial block. In the modified testbench, it was being set using a statement in the top-level generate block. # 04 - Verilog - Replacing a Constant with a Register (Verilog Basics) ## 04.1 - Summary ### Background: The first time the clock was toggled in this application, an output was toggled as expected, but it was followed by a 100ms delay. The second time the clock was toggled an output toggled as expected. The third time the clock was toggled, no output toggled. ### Initial Problem: The second time the clock toggled, the output toggled, but it was followed by a 100ms delay. ### Solution: The problem was caused by the testbench using a constant value for the delay. The value of the delay should have been a register because the register value is updated each time the clock is toggled. ## 04.2 - Code ### Verilog Code: module delay_test(input clk, output reg out); always @ (posedge clk) begin out<=~out; end endmodule ### Testbench Code: module delay_test(clk,out); reg clk, out; initial begin clk = 0; out = 0; end always begin #100 clk = ~clk; end endmodule ### Solution: The delay was due to the constant value being used for the delay. ### Solution: Instead of using a constant 100 for the delay, use a register and have the register value be updated each time the clock is toggled. ## 04.3 - Result ### Original: ### Modified: # 05 - Verilog - Creating a Sink - Writing a Testbench (Verilog Basics) ## 05.1 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Testbench Code: module sink_test(clk,out,in); reg clk, out, in; initial begin clk = 1; out = 4'b1111; in = 4'b0000; end always begin #100 clk = ~clk; in = in + 4'b0001; end endmodule ### Result: # 06 - Verilog - Creating a Sink - Writing a Functional Testbench (Verilog Basics) ## 06.1 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Functional Testbench Code: module sink_test(clk,out,in); reg clk, out, in; initial begin clk = 1; out = 4'b1111; in = 4'b0000; end always begin #100 clk = ~clk; in = in + 4'b0001; end initial begin $monitor(out = out, in = in); end initial $stop; endmodule ## 06.2 - Result: # 07 - Verilog - Creating a Sink - Reading a Functional Testbench (Verilog Basics) ## 07.1 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Functional Testbench Code: module sink_test(clk,out,in); reg clk, out, in; initial begin clk = 1; out = 4'b1111; in = 4'b0000; end always begin #100 clk = ~clk; in = in + 4'b0001; end initial begin $monitor(out = out, in = in); end initial $stop; endmodule ## 07.2 - Result: ## 07.3 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Functional Testbench Code: module sink_test(clk,out,in); reg clk, out, in; initial begin clk = 1; out = 4'b1111; in = 4'b0000; end always begin #100 clk = ~clk; in = in + 4'b0001; end initial begin $monitor(out = out, in = in); end initial $stop; endmodule ## 07.4 - Result: # 08 - Verilog - Creating a Sink - Reading a Testbench (Verilog Basics) ## 08.1 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Testbench Code: module sink_test(clk,out,in); reg clk, out, in; initial begin clk = 1; out = 4'b1111; in = 4'b0000; end always begin #100 clk = ~clk; in = in + 4'b0001; end initial begin $monitor(out = out, in = in); end initial $stop; endmodule ## 08.2 - Result: # 09 - Verilog - Creating Sinks in a Design Using a Module (Verilog Basics) ## 09.1 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Source Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end initial begin clk = 1; end always begin #100 clk = ~clk; in = in + 4'b0001; end initial begin $monitor(out = out, in = in); end initial $stop; endmodule ### Result: # 10 - Verilog - Creating Sinks in a Design Using a Module (Verilog Basics) ## 10.1 - Summary ### Verilog Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end always @ (posedge clk) begin out<=in; end endmodule ### Source Code: module sink_test(clk,out,in); reg [0:3] out; initial begin out = 4'b1111; end initial begin clk = 1; end always begin #100 clk = ~clk; in = in + 4'b0001; end initial begin $monitor(out = out, in = in); end initial $stop; endmodule ### Result: # 1