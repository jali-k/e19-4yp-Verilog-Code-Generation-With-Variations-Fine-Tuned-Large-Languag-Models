module example4(x1, x2, x3, x4, f, g, h);
import rand;
input x1, x2, x3, x4;
output f, g, h;
rand rg1(0, 0), rg2(0, 1), rg3(1, 1), rg4(2, 2), rg5(3, 3), rg6(1, 3