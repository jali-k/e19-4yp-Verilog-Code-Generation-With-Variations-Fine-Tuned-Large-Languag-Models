module gates4_top (
input wire [3:0] s1,
input wire [3:0] s2,
input wire [3:0] s3,
input wire [3:0] s4,
output wire [2:0] ld
);
gates4 U1
(
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0]),
.x()
);
wire[2:0] s = {s3, s4};
case(s1)
3'b0: s[0] = s1; break;
3'b1: s[0] = s2; break;
3'b2: s[0] = s3; break;
3'b3: s[0] = s4; break;
default: s[0] = s4; break;
endcase
case(s2)
3'b0: s[1] = s1; break;
3'b1: s[1] = s2; break;
3'b2: s[1] = s3; break;
3'b3: s[1] = s4; break;
default: s[1] = s4; break;
endcase
U2(
.x(s[0]),
.y(s[1]),
.and4_(ld[2]),
.or4_(ld[1]),
.xor4_(ld[0])
);
endmodule
### Execution Details:
The test bench, tb_gates4_top, is shown below. The input port is a 4 bit vector with two independent vectors from which to choose an operand. There are four cases, three of which involve using a constant, and the other using a constant index via an MDA.
When a constant is selected for operand, the test bench uses a constant index with a MDA to select the required operand.
When a constant index is selected for operand, the test bench uses an indexed port to indicate the operand.
### Execution Results:
The following results are generated by the test bench. For the first case, the constant index for operand is used. For the second case, the indexed port is used. In both cases, the same answer is generated which is correct.

## Summary:

If you can’t write and test a module, you aren’t a proper designer.

## References

[1] McLaren,.,, and. Digital Design with VHDL. Addison-Wesley, 2009.

[2]. Digital System Design: A Practical Approach Using VHDL and Verilog. Prentice Hall, 1999.

[3]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[4]  and. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[5]. VHDL tutorial. Addison-Wesley, 1993.

[6]. Digital Logic Design, 4th edition. Pearson, 2009.

[7]. A Handbook of VHDL Design, 2nd edition. Addison-Wesley, 2004.

[8] McLaren,.,, and. Digital Design with VHDL. Addison-Wesley, 2009.

[9]. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[10]. Digital Logic Design. Pearson, 1994.

[11]. Digital Design: A Practical Approach Using VHDL and Verilog. Prentice Hall, 1999.

[12]. Digital System Design: A Practical Approach Using VHDL and Verilog. Addison-Wesley, 2009.

[13]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[14]. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[15]. VHDL tutorial. Addison-Wesley, 1993.

[16]  and. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[17]. Digital Logic Design, 4th edition. Pearson, 2009.

[18]. A Handbook of VHDL Design, 2nd edition. Addison-Wesley, 2004.

[19]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[20]. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[21]. Digital Logic Design. Pearson, 1994.

[22]. Digital System Design: A Practical Approach Using VHDL and Verilog. Addison-Wesley, 2009.

[23]. VHDL tutorial. Addison-Wesley, 1993.

[24]  and. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[25]. Digital Logic Design, 4th edition. Pearson, 2009.

[26]. A Handbook of VHDL Design, 2nd edition. Addison-Wesley, 2004.

[27]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[28]. VHDL tutorial: a handbook.. Co., 1993.

[29]. Digital Logic Design. Pearson, 1994.

[30]. Digital System Design: A Practical Approach Using VHDL and Verilog. Addison-Wesley, 2009.

[31]. VHDL tutorial. Addison-Wesley, 1993.

[32]  and. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[33]. Digital Logic Design, 4th edition. Pearson, 2009.

[34]. A Handbook of VHDL Design, 2nd edition. Addison-Wesley, 2004.

[35]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[36]. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[37]. Digital Logic Design. Pearson, 1994.

[38]. Digital System Design: A Practical Approach Using VHDL and Verilog. Addison-Wesley, 2009.

[39]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[40]. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[41]. VHDL tutorial. Addison-Wesley, 1993.

[42]  and. VHDL tutorial: a handbook. Addison Wesley Pub. Co., 1993.

[43]. Digital Logic Design, 4th edition. Pearson, 2009.

[44]. A Handbook of VHDL Design, 2nd edition. Addison-Wesley, 2004.

[45]. VHDL, the very high level. New York: McGraw-Hill, 1989.

[46]. VHDL tutorial: a handbook.. Co., 1993.

[47]. Digital Logic Design. Pearson,