@gen_block1
module NOR5(