#### Testbench:
Test all the 32 combinatorial paths of the ALU4.
#### ALU4:
Test all the 32 combinatorial paths of the ALU4.