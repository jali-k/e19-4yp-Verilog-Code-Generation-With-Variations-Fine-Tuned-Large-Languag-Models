```verilog
module aoi2(g,a,b,c,d,e);
output g;
input a,b,c,d;
wire [0:3] e;

// Dataflow assignments for