The modified code can be found in the `Modified` branch.