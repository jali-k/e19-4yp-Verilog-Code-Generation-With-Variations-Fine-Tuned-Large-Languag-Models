enum {off, on} state;

Reset_Prog M1 (clk, resetn, state);
### Result
**
```
### [Top](#top)
### [Next](#next)
### [Next](#next)
### [Next](#next)
### [Next](#next)
### [Next](#next)
### [Next](#next)
### [Next](#next)