{% include_relative cmp.v %}
### Testbench Code:
{% include_relative tb_TOP1.v %}
### Input Log:
{% include_relative cmp.log %}
### Output Log:
{% include_relative cmp.out %}
### Expected Result:
* 0: 1
* 1: 0
* 2: 0
* 3: 1
* 4: 1
* 5: 1
* 6: 1
* 7: 1
* 8: 1
* 9: 0