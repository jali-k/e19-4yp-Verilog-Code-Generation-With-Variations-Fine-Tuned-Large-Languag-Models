module DataComponent (Data