initial begin