module example7_13(D