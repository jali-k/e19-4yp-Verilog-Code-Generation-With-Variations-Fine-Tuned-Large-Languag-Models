```
module show_aa(ao,ai); // NOT gate with delay 2
  output ao; input ao;
  show_aa ao,ai;
endmodule
```
### Test Inputs:
![image](https://user-images.githubusercontent.com/62660481/215289069-7d9ec12d-c37a-45a5-8f3c-d68b0fc2e918.png)