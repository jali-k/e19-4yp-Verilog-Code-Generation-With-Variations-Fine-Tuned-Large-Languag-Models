int func(int f, int x3, int x2, int x1)
{
    if ((x2 == 0) && (x1 == 1)) {
	f = x3;
    } else {
	f =