module Xoring (input a, b, output y);