module test_k;
wire q, clock, j, k, preset, clear;
reg j, k;
jkEdge