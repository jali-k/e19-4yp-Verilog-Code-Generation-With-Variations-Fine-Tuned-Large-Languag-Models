if(i2 == a [j+:3]) // Added inside
### Modified Simulation:
$readmemb("test_vector.txt",a);
j=1; // Added
i2=a[j+:3];
$monitor($time,"i1=%b,i2=%b,o=%b",i1,i2,o);
Initialization:
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i1=0;
i2=0;
i