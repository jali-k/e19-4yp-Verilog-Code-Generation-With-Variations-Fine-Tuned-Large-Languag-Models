```verilog
`timescale 1ns/100ps
module Comparator (input logic CLK, RST_X,