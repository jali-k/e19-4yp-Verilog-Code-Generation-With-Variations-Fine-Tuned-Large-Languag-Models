interface intf(input logic clk);
  logic s, ca;
endinterface

module tstha_9(intf.in intf1, input data);
  ha_