```Verilog
module wire_assign( input bit reset, input bit clk, output bit out