`module gade(a,a1,b,c,b1,c1);
interface iface();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface1();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface2();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface3();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface4();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface5();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface6();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface7();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface8();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface9();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface10();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface11();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface12();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface13();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface14();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface15();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface16();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface17();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface18();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface19();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface20();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface21();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface22();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface23();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface24();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface25();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface26();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface27();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface28();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface29();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface30();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface31();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface32();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface33();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface34();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface35();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface36();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface37();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface38();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface39();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface40();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface41();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface42();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface43();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface44();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface45();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface46();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface47();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface48();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface49();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface50();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface51();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface52();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface53();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface54();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface55();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface56();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface57();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface58();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface59();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface60();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface61();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface62();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface63();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface64();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface65();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface66();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface67();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface68();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface69();
logic b,c,b1,c1;
logic a,a1;
endinterface
interface iface70();
logic