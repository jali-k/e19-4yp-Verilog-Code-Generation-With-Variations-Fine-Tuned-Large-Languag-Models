module mux4to1(w0, w1, w2, w3, S, f);
input w0, w1, w2, w3;
input [1:0] S;
output f;
reg f;
localparam packed [1:0] selects = {2'b00, 2'b01, 2'b10, 2'b11};
always @(w0 or w1 or w2 or w3 or S)
    f = inside(S, selects);
endmodule