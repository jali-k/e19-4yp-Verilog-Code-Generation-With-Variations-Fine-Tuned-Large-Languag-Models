module testbench ();
generate data;
struct { rand int rand_member; } t1;
process data;
endmodule