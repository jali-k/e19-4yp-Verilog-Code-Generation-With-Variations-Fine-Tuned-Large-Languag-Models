module testbench ();
struct { rand bit[7:0] value;  } data;
process data;