module mux21b (
input wire a,
input wire b,
input wire s,
output reg y // Output must be reg for procedural assignment
);
always @(*) // Combinational sensitivity
case(s)
0: y = a; // Select a if s=0
1: y = b; // Select b if s=1
endcase
endmodule
### Results:
1. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux is set to 0 and 1.
2. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
3. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
4. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
5. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
6. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
7. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
8. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
9. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
10. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
11. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
12. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
13. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
14. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
15. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
16. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
17. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
18. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
19. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
20. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
21. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
22. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
23. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
24. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
25. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
26. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
27. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
28. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the 21mux of course being 3 in both cases.
29. 
The simulation tool was used to generate a waveform on the output port of a 32x32 21mux. The outputs of the 21mux are set to 0 and 1 along with the address line of the