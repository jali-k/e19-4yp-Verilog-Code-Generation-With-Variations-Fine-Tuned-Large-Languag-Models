`generate` for i in 0 to 15 generate s_