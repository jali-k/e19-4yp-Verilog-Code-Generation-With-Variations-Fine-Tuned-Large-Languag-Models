module dff_with_reset(data, clock, r, out);
input clock, r, data;
output out;
reg out;
always @(posedge clock or posedge r)
begin
if (r)
out = 0;
else if(data inside {1, [1]})
out = data;
end
endmodule
### Output:
0001 1111 1010 1001 1101 1100 0100 0100 0010 1111 1101 1010 0011 1101 0010 1101 0100 1111 1011 0011 
0001 1111 1010 1001 1101 1100 0100 0100 0010 1111 1101 1010 0011 1101 0010 1101 0100 1111 1011 0011 
### Generated by VERDI