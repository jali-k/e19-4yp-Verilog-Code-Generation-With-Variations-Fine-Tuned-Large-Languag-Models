${C_VAR,"<?=`C_VAR`?>".substr(1).escaped}.(a,clk,N, En) ${C_VAR,"<?=`C_VAR`?>".substr(C_VAR.size-1).escaped, C_VAR}.(<?, a, [N : 0]>,clk, En);
### Simulation Results:
### Logic Synthesis Results:
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
### 
###