module Clock_Mod_12();
initial
begin
name_b: