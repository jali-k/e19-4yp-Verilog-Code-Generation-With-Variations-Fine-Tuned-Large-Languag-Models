// DFF with async preset
module dffalter_tst(); // Testbench, likely for a DFF named dffalter
reg di,clk,clr,pr;
wire q, qb; // Added qb
// dffalter dff(q,qb,di,clk,clr,pr); // Assumed instantiation of DUT
initial
begin
clr=1'b1;pr=1'b0;clk=1'b0;di=1'b0; // Start with clear asserted
end
always
begin
clr=1'b0; // Deassert clear
end
always #16 pr=1'b1; // Assert preset
always #20 pr =1'b0; // Deassert preset
always # 4 di =~di; // Toggle data
initial $monitor("t=%0d, clk=%b, clr=%b, pr=%b, di=%b, q=%b ", $time,clk,clr,pr,di,q);
initial #46 $stop; // Stop simulation
endmodule
### Inserted Code:
// Async preset behavior
module dffalter_tst(); // Testbench, likely for a DFF named dffalter
reg di,clk,clr,pr;
wire q, qb; // Added qb
// dffalter dff(q,qb,di,clk,clr,pr); // Assumed instantiation of DUT
initial
begin
clr=1'b1;pr=1'b0;clk=1'b0;di=1'b0; // Start with clear asserted
end
always
begin
clr=1'b0; // Deassert clear
end
always # 4 di =~di; // Toggle data
always #16 pr=1'b1; // Assert preset
always #20 pr =1'b0; // Deassert preset
initial $monitor("t=%0d, clk=%b, clr=%b, pr=%b, di=%b, q=%b pkg.di=%b ", $time,clk,cl