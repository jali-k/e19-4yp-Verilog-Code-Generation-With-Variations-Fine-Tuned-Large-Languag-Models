module dff_inst(D, Clock, Resetn, Q);
input D, Clock, Resetn;
output Q