module Sched