module ALU (output[31:0] Result, input[31:0] ArgA, ArgB, input Clk);
specify
    specparam tRise = 9, tFall = 4;
    (Clk *> Result) = (tRise, tFall);
    signed [3:0] a, b;
    logic[3:0] b1, b2, b3, b4;
    a = ArgA[31:0];
    b = ArgB[31:0];
    assign {b3, b2, b1, b4} = ArgA[3:0];
    assign {b[3], b[2], b[1], b[0]} = b2;
    assign {b[3], b[2], b[1], b[0]} = b1;
    assign {b3, b2, b1, b4} = b4;
    (a(3), a(2), a(1), a(0)) = b2[3:0];
    (b(3), b(2), b(1), b(0)) = b1[3:0];
    logic [2:0] b5, b6, b7;
    assign {b5, b6, b7} = ArgB[3:0];
    assign b6 = ArgB[0];
    assign b7 = ArgB[1];
endspecify
endmodule

```

The following are the results.

```
# 1059001_1.v
# 1059002_1.v
# 1059003_1.v
#
# 1059001_2.v
# 1059002_2.v
# 1059003_2.v
#
# 1059001_3.v
# 1059002_3.v
# 1059003_3.v
#
# 1059001_4.v
# 1059002_4.v
# 1059003_4.v
#
# 1059001_5.v
# 1059002_5.v
# 1059003_5.v
#
# 1059001_6.v
# 1059002_6.v
# 1059003_6.v
#
# 1059001_7.v
# 1059002_7.v
# 1059003_7.v
#
# 1059001_8.v
# 1059002_8.v
# 1059003_8.v
#
# 1059001_9.v
# 1059002_9.v
# 1059003_9.v
#
# 1059001_10.v
# 1059002_10.v
# 1059003_10.v
#
# 1059001_11.v
# 1059002_11.v
# 1059003_11.v
#
# 1059001_12.v
# 1059002_12.v
# 1059003_12.v
#
# 1059001_13.v
# 1059002_13.v
# 1059003_13.v
#
# 1059001_14.v
# 1059002_14.v
# 1059003_14.v
#
# 1059001_15.v
# 1059002_15.v
# 1059003_15.v
#
# 1059001_16.v
# 1059002_16.v
# 1059003_16.v
#
# 1059001_17.v
# 1059002_17.v
# 1059003_17.v
#
# 1059001_18.v
# 1059002_18.v
# 1059003_18.v
#
# 1059001_19.v
# 1059002_19.v
# 1059003_19.v
#
# 1059001_20.v
# 1059002_20.v
# 1059003_20.v
#
# 1059001_21.v
# 1059002_21.v
# 1059003_21.v
#
# 1059001_22.v
# 1059002_22.v
# 1059003_22.v
#
# 1059001_23.v
# 1059002_23.v
# 1059003_23.v
#
# 1059001_24.v
# 1059002_24.v
# 1059003_24.v
#
# 1059001_25.v
# 1059002_25.v
# 1059003_25.v
#
# 1059001_26.v
# 1059002_26.v
# 1059003_26.v
#
# 1059001_27.v
# 1059002_27.v
# 1059003_27.v
#
# 1059001_28.v
# 1059002_28.v
# 1059003_28.v
#
# 1059001_29.v
# 1059002_29.v
# 1059003_29.v
#
# 1059001_30.v
# 1059002_30.v
# 1059003_30.v
#
# 1059001_31.v
# 1059002_31.v
# 1059003_31.v
#
# 1059001_32.v
# 1059002_32.v
# 1059003_32.v
#
# 1059001_33.v
# 1059002_33.v
# 1059003_33.v
#
# 1059001_34.v
# 1059002_34.v
# 1059003_34.v
#
# 1059001_35.v
# 1059002_35.v
# 1059003_35.v
#
# 1059001_36.v
# 1059002_36.v
# 1059003_36.v
#
# 1059001_37.v
# 1059002_37.v
# 1059003_37.v
#
# 10