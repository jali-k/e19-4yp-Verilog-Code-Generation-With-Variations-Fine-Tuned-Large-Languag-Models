// Verilog code for Problem 11
module Full_Subtractor(
    input logic A