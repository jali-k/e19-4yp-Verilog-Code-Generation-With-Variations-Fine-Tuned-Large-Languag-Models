always @( posedge clk ) begin : clocked
deassign