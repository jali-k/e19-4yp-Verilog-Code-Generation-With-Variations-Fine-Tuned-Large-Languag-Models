```v
module TOP1(CLK, RST_X);
  // Inputs
  input CLK;
  input RST_X;

  // Outputs
  // Verilog Code Generation

  // Verilog Code Generation
  // Instantiate the verilog code to be included in the module definition

  // Parameters

  // Localparam

  // Variables

  // Direct memories

  // Generated code

  localparam TOP1_x_array_0 = 1;

  localparam TOP1_x_array_1 = 2;

  localparam TOP1_x_array_2 = 3;

  localparam TOP1_x_array_3 = 4;

  localparam TOP1_x_array_4 = 5;

  localparam TOP1_x_array_5 = 6;

  localparam TOP1_x_array_6 = 7;

  localparam TOP1_x_array_7 = 8;

  localparam TOP1_x_array_8 = 9;

  localparam TOP1_x_array_9 = 10;

  localparam TOP1_x_array_10 = 11;

  localparam TOP1_x_array_11 = 12;

  localparam TOP1_x_array_12 = 13;

  localparam TOP1_x_array_13 = 14;

  localparam TOP1_x_array_14 = 15;

  localparam TOP1_x_array_15 = 16;

  localparam TOP1_x_array_16 = 17;

  localparam TOP1_x_array_17 = 18;

  localparam TOP1_x_array_18 = 19;

  localparam TOP1_x_array_19 = 20;

  localparam TOP1_x_array_20 = 21;

  localparam TOP1_x_array_21 = 22;

  localparam TOP1_x_array_22 = 23;

  localparam TOP1_x_array_23 = 24;

  localparam TOP1_x_array_24 = 25;

  localparam TOP1_x_array_25 = 26;

  localparam TOP1_x_array_26 = 27;

  localparam TOP1_x_array_27 = 28;

  localparam TOP1_x_array_28 = 29;

  localparam TOP1_x_array_29 = 30;

  localparam TOP1_x_array_30 = 31;

  localparam TOP1_x_array_31 = 32;

  localparam TOP1_x_array_32 = 33;

  localparam TOP1_x_array_33 = 34;

  localparam TOP1_x_array_34 = 35;

  localparam TOP1_x_array_35 = 36;

  localparam TOP1_x_array_36 = 37;

  localparam TOP1_x_array_37 = 38;

  localparam TOP1_x_array_38 = 39;

  localparam TOP1_x_array_39 = 40;

  localparam TOP1_x_array_40 = 41;

  localparam TOP1_x_array_41 = 42;

  localparam TOP1_x_array_42 = 43;

  localparam TOP1_x_array_43 = 44;

  localparam TOP1_x_array_44 = 45;

  localparam TOP1_x_array_45 = 46;

  localparam TOP1_x_array_46 = 47;

  localparam TOP1_x_array_47 = 48;

  localparam TOP1_x_array_48 = 49;

  localparam TOP1_x_array_49 = 50;

  localparam TOP1_x_array_50 = 51;

  localparam TOP1_x_array_51 = 52;

  localparam TOP1_x_array_52 = 53;

  localparam TOP1_x_array_53 = 54;

  localparam TOP1_x_array_54 = 55;

  localparam TOP1_x_array_55 = 56;

  localparam TOP1_x_array_56 = 57;

  localparam TOP1_x_array_57 = 58;

  localparam TOP1_x_array_58 = 59;

  localparam TOP1_x_array_59 = 60;

  localparam TOP1_x_array_60 = 61;

  localparam TOP1_x_array_61 = 62;

  localparam TOP1_x_array_62 = 63;

  localparam TOP1_x_array_63 = 64;

  localparam TOP1_x_array_64 = 65;

  localparam TOP1_x_array_65 = 66;

  localparam TOP1_x_array_66 = 67;

  localparam TOP1_x_array_67 = 68;

  localparam TOP1_x_array_68 = 69;

  localparam TOP1_x_array_69 = 70;

  localparam TOP1_x_array_70 = 71;

  localparam TOP1_x_array_71 = 72;

  localparam TOP1_x_array_72 = 73;

  localparam TOP1_x_array_73 = 74;

  localparam TOP1_x_array_74 = 75;

  localparam TOP1_x_array_75 = 76;

  localparam TOP1_x_array_76 = 77;

  localparam TOP1_x_array_77 = 78;

  localparam TOP1_x_array_78 = 79;

  localparam TOP1_x_array_79 = 80;

  localparam TOP1_x_array_80 = 81;

  localparam TOP1_x_array_81 = 82;

  localparam TOP1_x_array_82 = 83;

  localparam TOP1_x_array_83 = 84;

  localparam TOP1_x_array_84 = 85;

  localparam TOP1_x_array_85 = 86;

  localparam TOP1_x_array_86 = 87;

  localparam TOP1_x_array_87 = 88;

  localparam TOP1_x_array_88 = 89;

  localparam TOP1_x_array_89 = 90;

  localparam TOP1_x_array_90 = 91;

  localparam TOP1_x_array_91 = 92;

  localparam TOP1_x_array_92 = 93;

  localparam TOP1_x_array_93 = 94;

  localparam TOP1_x_array_94 = 95;

  localparam TOP1_x_array_95 = 96;

  localparam TOP1_x_array_96 = 97;

  localparam TOP1_x_array_97 = 98;

  localparam TOP1_x_array_98 = 99;

  localparam TOP1_x_array_99 = 100;

  localparam TOP1_x_array_100 = 101;

  localparam TOP1_x_array_101 = 102;

  localparam TOP1_x_array_102 = 103;

  localparam TOP1_x_array_103 = 104;

  localparam TOP1_x_array_104 = 105;

  localparam TOP1_x_array_105 = 106;

  localparam TOP1_x_array_106 = 107;

  localparam TOP1_x_array_107 = 108;

  localparam TOP1_x_array_108 = 109;

  localparam TOP1_x_array_109 = 110;

  localparam TOP1_x_array_110 = 111;

  localparam TOP1_x_array_111 = 112;

  localparam TOP1_x_array_112 = 113;

  localparam TOP1_x_array_113 = 114;

  localparam TOP1_x_array_114 = 115;

  localparam TOP1