// Create a module with one input and one output that behaves like a wire
module wire_assign_bit( input in, output out );
    // assign out to in
    assign out = in;
endmodule
/Lab/Lab2_Arijit/Lab2_Arijit/testbench.h
//
//  testbench.h
//  Lab2_Arijit
//
//  Created by  on 11/19/14.
//  Copyright (c) 2014. All rights reserved.
//

#ifndef __Lab2_Arijit__testbench__
#define __Lab2_Arijit__testbench__

#include <iostream>

#endif /* defined(__Lab2_Arijit__testbench__) */