module reg8(D, Clock, Resetn, Q);
input [