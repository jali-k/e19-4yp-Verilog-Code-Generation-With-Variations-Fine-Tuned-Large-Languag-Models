```Verilog
module shift_reg( input [3:0] d_in, input clk