module fulladder(a,b,c,s,carry);
input a,b