module adder4(
input wire a,
input wire b,
input wire ci,
input