module example5(x1, x2, x3, f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
    if (x2 == 1)
        f = x1;
    else if (x2 >= 2 && x2 <= 3)
        f = x3;
    end
endmodule
### New Code:
module example5(x1, x2, x3, f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
    if (x2 >= 2 && x2 <= 3)
        f = x3;
    else if (x2 == 1)
        f = x1;
    end
endmodule
### End Time: 07:46
"""

# TODO: Implement the solution logic here.
# This dictionary should contain the final modified code for each example.
# The key to this dictionary should be the title of the test case.
# The value should be the string of the modified code.
solution = {}
"""
#This code is generated using the Variation: Add an if block testing whether part-select of a packed array is inside a fixed constant range.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 >= 2 && x2 <= 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 1 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 2 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 == 2)
f = x2;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 3 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 == 2)
f = x2;
else if (x2 == 3)
f = x3;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 4 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 == 2)
f = x2;
else if (x2 == 3)
f = x3;
else if (x2 == 4)
f = x4;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
"""
solution['example5'] = """
#This code is generated using the Variation: Add an if block testing whether part-select of a packed array is inside a fixed constant range.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 >= 2 && x2 <= 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 1 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 2 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 == 2)
f = x2;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 3 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 == 2)
f = x2;
else if (x2 == 3)
f = x3;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
    #This code is generated using the Variation: Add a new test case with only one input signal of 4 and no other signals.
#The Original code is:
module example5(x1, x2, x3,
f);
input x1, x2, x3;
output f;
reg f;
always @(x1 or x2 or x3)
if (x2 == 1)
f = x1;
else if (x2 == 2)
f = x2;
else if (x2 == 3)
f = x3;
else if (x2 == 4)
f = x4;
else if (x2 < 2 && x2 > 3)
f = x3;
end
endmodule
"""

# Save your solution:
solution_path = "assignment7_solution.py"

with open(solution_path, "w") as solution_file:
    solution_file.write("# DO NOT MODIFY THIS FILE\n")
    solution_file.write("# This file was automatically generated by assignment7.py\n")
    solution_file.write("solution = {}\n".format(solution))

print("Solution written to {}".format(solution_path))
print("Please add this file to your git repo.  You can do this in two steps.")
print("Step 1: go to the directory containing this file and run")
print("    git add {}".format(solution_path))
print("Step 2: go to your github.com repository and click 'Create Pull Request'")
#!git add assignment7_solution.py

#!git commit -m "assignment7_solution.py, final"

#!git push

# + [markdown] nbgrader={"grade": false, "locked": true, "solution": false}
# ## Submission Instructions
#
# Make sure you fill in any place that says `YOUR CODE HERE` or "YOUR ANSWER HERE", as well as your name and collaborators below:

# + nbgrader={"grade": false, "locked": false, "solution": false}
YOUR_ID = "00000000" # please fill here YOUR_ID
YOUR_COLLABORATORS =