`module Multiplier4 (input [1:0] A, B, input [7:0] Cin, output reg [3:0] Result, output reg CarryOut);
input [7:0] X, Y, Cin;
reg [31:0] Sum;