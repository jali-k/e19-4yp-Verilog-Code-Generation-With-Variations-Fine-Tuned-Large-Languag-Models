module hex7seg_le (
input wire [3:0] x,
output wire [6:0] a_to_g // Outputs for segments a,b,c,d,e,f,g
);
genvar i;
generate
for(i=0; i<4; i++) :
begin: inside
assign a_to_g[6] = x[i] & ~x[3-i]; // a (segment index 6)
end
endgenerate
assign a_to_g[5] = x[2] & x[1] & ~x[0] // b (segment index 5)
| x[3] & x[1] & x[0]
| ~x[3] & x[2] & ~x[1] & x[0]
| x[3] & x[2] & ~x[1] & ~x[0];
assign a_to_g[4] = ~x[3] & ~x[2] & x[1] & ~x[0] // c (segment index 4)
| x[3] & x[2] & x[1]
| x[3] & x[2] & ~x[0];
assign a_to_g[3] = ~x[3] & ~x[2] & ~x[1] & x[0] // d (segment index 3)
| ~x[3] & x[2] & ~x[1] & ~x[0]
| x[3] & ~x[2] & x[1] & ~x[0]
| x[2] & x[1] & x[0];
assign a_to_g[2] = ~x[3] & x[0] // e (segment index 2)
| ~x[3] & x[2] & ~x[1]
| ~x[2] & ~x[1] & x[0];
assign a_to_g[1] = ~x[3] & ~x[2] & x[0] // f (segment index 1)
| ~x[3] & ~x[2] & x[1]
| ~x[3] & x[1] & x[0]
| x[3] & x[2] & ~x[1] & x[0];
assign a_to_g[0] = ~x[3] & ~x[2] & ~x[1] // g (segment index 0)
| x[3] & x[2] & ~x[1] & ~x[0]
| ~x[3] & x[2] & x[1] & x[0];
endmodule