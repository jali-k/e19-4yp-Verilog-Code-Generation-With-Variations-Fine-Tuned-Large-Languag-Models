module xor(out,a,b); // module for XOR gate
  input a,b;
  output out;
  xor a b out;
  endmodule
### Results:
<center>
<img src="img/11.png" width="500"