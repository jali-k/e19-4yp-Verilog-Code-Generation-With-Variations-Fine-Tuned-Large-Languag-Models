module add