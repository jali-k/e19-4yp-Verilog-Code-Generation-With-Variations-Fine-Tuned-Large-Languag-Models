```vhdl