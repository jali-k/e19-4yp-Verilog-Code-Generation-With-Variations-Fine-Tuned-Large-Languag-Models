```verilog
module nil;
reg [1:0]