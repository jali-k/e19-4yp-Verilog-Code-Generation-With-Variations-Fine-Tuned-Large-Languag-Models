[Verilog Code](anding_union_packed.v)

### Simulation:
![anding_union_packed](./images/anding_union_packed.png)

### Test Suite:
[Test Suite](anding_union_packed_testbench_suite.v)




## 4 Summary

In this Tutorial you have learned to use the following:

- Union
- Packed Union
- Use packed union as module port
- Use packed union as module input

Note that these concepts can be used in the same manner in Verilog and VHDL.

## 5 References

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=176&zoom=auto,-230,1001)

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=176&zoom=auto,-230,1001)

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=176&zoom=auto,-230,1001)

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=176&zoom=auto,-230,1001)

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=176&zoom=auto,-230,1001)

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=176&zoom=auto,-230,1001)

[Xilinx - Verilog Union](https://www.xilinx.com/support/documentation/user_guides/ug478_7Series_Config.pdf#page=17