module net_gate(x,y,z);
input x,y;
output [2:1] z;
wire [1:0] nn;
and (nn,x,y);
assign z=nn[0];
endmodule
### Result:
Error: net_gate.v(13) : syntax error, unexpected IDENT([2:1]), expecting {identifier(104), (identifier(104), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (constant_any(175), (, identifier(104), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, constant_any(175), (, ), identifier(104), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175)), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant_any(175), (, ), constant