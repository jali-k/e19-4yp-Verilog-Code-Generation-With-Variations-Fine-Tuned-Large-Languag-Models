module JerkyComparator(output[1:0] AdjustFreq, input ClockIn, PLLClock, Reset);
reg[1:0] Adjr;
assign AdjustFreq = Adjr;
reg[1:0] HiCount;
always @(ClockIn, Reset)
if (Reset==1'b1)
begin
    Adjr = 2'b01;
    HiCount = 2'b0;
end
else if (PLLClock==1'b1)
    HiCount = HiCount + 2'b01;
else begin
    case (HiCount)
        2'b00: Adjr = 2'b11;
        2'b01: Adjr = 2'b01;
        default: Adjr = 2'b00;
    endcase
    HiCount = 2'b0;
end
endmodule
#100000001
#100000002
#100000003
#100000004
#100000005
#100000006
#100000007
#100000008
#100000009
#100000010
#100000011
#100000012
#100000013
#100000014
#100000015
#100000016
#100000017
#100000018
#100000019
#100000020
#100000021
#100000022
#100000023
#100000024
#100000025
#100000026
#100000027
#100000028
#100000029
#100000030
#100000031
#100000032
#100000033
#100000034
#100000035
#100000036
#100000037
#100000038
#100000039
#100000040
#100000041
#100000042
#100000043
#100000044
#100000045
#100000046
#100000047
#100000048
#100000049
#100000050
#100000051
#100000052
#100000053
#100000054
#100000055
#100000056
#100000057
#100000058
#100000059
#100000060
#100000061
#100000062
#100000063
#100000064
#100000065
#100000066
#100000067
#100000068
#100000069
#100000070
#100000071
#100000072
#100000073
#100000074
#100000075
#100000076
#100000077
#100000078
#100000079
#100000080
#100000081
#100000082
#100000083
#100000084
#100000085
#100000086
#100000087
#100000088
#100000089
#100000090
#100000091
#100000092
#100000093
#100000094
#100000095
#100000096
#100000097
#100000098
#100000099
#100000100
#100000101
#100000102
#100000103
#100000104
#100000105
#100000106
#100000107
#100000108
#100000109
#100000110
#100000111
#100000112
#100000113
#100000114
#100000115
#100000116
#100000117
#100000118
#100000119
#100000120
#100000121
#100000122
#100000123
#100000124
#100000125
#100000126
#100000127
#100000128
#100000129
#100000130
#100000131
#100000132
#100000133
#100000134
#100000135
#100000136
#100000137
#100000138
#100000139
#100000140
#100000141
#100000142
#100000143
#100000144
#100000145
#100000146
#100000147
#100000148
#100000149
#100000150
#100000151
#100000152
#100000153
#100000154
#100000155
#100000156
#100000157
#100000158
#100000159
#100000160
#100000161
#100000162
#100000163
#100000164
#100000165
#100000166
#100000167
#100000168
#10