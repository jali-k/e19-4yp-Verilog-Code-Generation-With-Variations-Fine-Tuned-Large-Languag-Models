// Verilog code for Problem 5
module Half