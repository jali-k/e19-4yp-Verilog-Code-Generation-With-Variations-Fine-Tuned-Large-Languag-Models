module XOR1(out,in1,in2);