module func1(x1, x2, x3, f);
input x1, x2, x3