```verilog
module full_adder(i1, i2, cin, sum, cout);
input i1, i2