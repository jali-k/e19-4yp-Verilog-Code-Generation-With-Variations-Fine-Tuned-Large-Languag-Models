module testbench ();
generate struct { rand bit [3:0] fork statement;} fork statement;
process fork statement;
endmodule
### Base Verilog Code:
module testbench ();
generate fork join_any