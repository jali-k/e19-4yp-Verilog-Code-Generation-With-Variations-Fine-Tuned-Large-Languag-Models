module dffalter_tst(in wire clk, inout wire q, inout wire qb, in out wire di, in out wire clr, in out wire pr);
import mypkg::*;
reg qb,q;
assign qb=q[1:0];
assign q[1:0]=di[1:0];
// dffalter dff(q,qb,di,clk,clr,pr);
initial
begin
clr=1'b0;pr=1'b0; // Start with preset and clear deasserted
end
always
begin
clr=1'b0; // Deassert clear
end
always # 4 di =~di; // Toggle data
always #16 pr=1'b1; // Assert preset
always #20 pr =1'b0; // Deassert preset
initial
begin
$monitor("**t=%0d, clk=%b, clr=%b, pr=%b, di=%b, q=%b, qb=%b ", $time,clk,clr,pr,di[1:0],q[1:0],qb[1:0]);
end
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");
initial $monitor("**");