module test_carry;
reg a, b, c;
integer i;
wire cout;
generate
carry c1(cout, c, a, b);
endgenerate
endmodule
### Result:
**Time** : 0 ns
**Output:**
**a** : x
**b** : x
**c** : 0
**cout** : 0
**a** : x
**b** : x
**c** : 0
**cout** : 0
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 0
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** : 1
**b** : 1
**c** : 1
**cout** : 1
**a** :