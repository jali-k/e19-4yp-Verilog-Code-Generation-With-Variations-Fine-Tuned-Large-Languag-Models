module tst_nm_in();
  reg in; wire out;

  parameter NUM_P = 16;
  parameter NUM_N = 16;

  reg [NUM_P-1:0] P[NUM_N-1:0];
  reg [NUM_N-1:0] N[NUM_P-1:0];

  reg [NUM_P-1:0] Q;
  reg [NUM_N-1:0] R;

  wire [NUM_P-1:0] S_NM;
  wire [NUM_N-1:0] X_NM;

  wire [NUM_P-1:0] S_PN;
  wire [NUM_N-1:0] X_PN;

  wire [NUM_P-1:0] S_NN;
  wire [NUM_N-1:0] X_NN;

  reg [NUM_P-1:0] S_NM_P;
  wire [NUM_N-1:0] X_NM_P;

  reg [NUM_P-1:0] S_PN_P;
  wire [NUM_N-1:0] X_PN_P;

  wire [NUM_P-1:0] S_NN_P;
  wire [NUM_N-1:0] X_NN_P;

  wire [NUM_P-1:0] S_NM_N;
  wire [NUM_N-1:0] X_NM_N;

  wire [NUM_P-1:0] S_PN_N;
  wire [NUM_N-1:0] X_PN_N;

  wire [NUM_P-1:0] S_NN_N;
  wire [NUM_N-1:0] X_NN_N;

  NMOSinv_1 nmv1(
    X_NM,
    in,
    S_NM,
    NUM_P,
    NUM_N,
    P,
    N,
    Q,
    NUM_N,
    X_NM_N,
    NUM_P,
    X_NM_P,
    NUM_P,
    S_NM_N,
    X_PN_P,
    S_NM_P,
    Q,
    X_PN,
    NUM_N,
    NUM_P,
    NUM_N,
    X_NN_N,
    X_PN_N,
    X_NN_P);

  NMOSinv_1 nmv2(
    X_NN,
    NUM_N,
    NUM_P,
    X_NN_N,
    NUM_N,
    S_NN,
    NUM_P,
    X_NN_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_P,
    NUM_N,
    P,
    NUM_P,
    NUM_N,
    X_PN_N,
    Q,
    S_PN,
    NUM_P,
    X_PN,
    NUM_N,
    NUM_N,
    X_NM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    X_NM_P,
    NUM_P,
    X_NM,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    P,
    X_PN_P,
    X_NM_N,
    NUM_P,
    NUM_N,
    S_PN_P,
    S_NM_N,
    X_PN_N,
    S_PN_N,
    S_PN_N,
    S_PN_N,
    X_NN_P,
    X_NN_N,
    X_NN_N,
    X_NN_N,
    S_NM_N);

  NMOSinv_1 nmv3(
    X_NM_P,
    NUM_P,
    NUM_N,
    X_NM_N,
    S_NM_N,
    X_PN_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    P,
    NUM_P,
    S_NM_P,
    Q,
    NUM_N,
    S_PN_P,
    NUM_N,
    N,
    X_NN_N,
    X_PN_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    X_NN_P,
    X_NN_N,
    NUM_N,
    NUM_P,
    NUM_P,
    X_PN_P,
    X_NM_N,
    NUM_P,
    NUM_N);

  NMOSinv_1 nmv4(
    X_PN,
    NUM_N,
    NUM_P,
    X_PN_N,
    NUM_N,
    X_NN_N,
    NUM_P,
    NUM_P,
    NUM_P,
    NUM_N,
    S_PN,
    NUM_N,
    X_PN_P,
    X_NN_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    X_NN_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_P,
    NUM_N);

  NMOSinv_1 nmv5(
    X_NN_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    X_PN_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_P);

  NMOSinv_1 nmv6(
    S_PN_P,
    NUM_P,
    NUM_N,
    X_PN_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    X_PN_P,
    NUM_P,
    NUM_N,
    X_PN_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    S_PN_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_P);

  NMOSinv_1 nmv7(
    S_NN_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_P);

  NMOSinv_1 nmv8(
    X_NM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_N,
    NUM_P,
    NUM_P,
    NUM_P,
    NUM_N,
    NUM_P,
    NUM_N);

  NMOSinv_1 nmv9(
    F2_S(
      NUM_P,
      NUM_N,
      P,
      NUM_N,
      S_PN,
      NUM_N,
      N,
      NUM_P,
      NUM_P,
      X_NN_N,
      NUM_N,
      S_NN,
      Q,
      NUM_N,
      X_PN_N,
      NUM_N,
      NUM_N,
      NUM_N,
      NUM_P,
      NUM_N,
      NUM_P,
      NUM_P,
      NUM_P,
      NUM_P,
      NUM_N,
      NUM_N,
      NUM_P,
      NUM_P,
      NUM_N,
      NUM_P,
      NUM_N,
      NUM_N,
      NUM_P,
      NUM_P,
      NUM_P,
      NUM_N,
      NUM_N