module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;// a1,a2,b1,b2 form the input
//ports of the module
output o;//o is the single output port of the module
wire o1,o2;//o1 and o2 are intermediate signals
//within the module
and g1(o1,a1,a2); //The AND gate primitive has two
and g2(o2,b1,b2);// instantiations with assigned
//names g1 & g2.
nor g3(o,o1,o2);//The nor gate has one instantiation
//with assigned name g3.
endmodule
### Verified Code:
module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;
output o;
wire o1,o2;
and g1(o1,a1,a2);
and g2(o2,b1,b2);
nor g3(o,o1,o2);
endmodule
### Violated Code:
module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;
output o;
wire o1,o2;
and g1(o1,a1,a2);
and g2(o2,b1,b2);
nor g3(o,o1,o2);
endmodule
### Violated Code:
module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;
output o;
wire o1,o2;
and g1(o1,a1,a2);
and g2(o2,b1,b2);
nor g3(o,o1,o2);
endmodule
### Violated Code:
module aoi_gate(o,a1,a2,b1,b2);
input a1,a2,b1,b2;
output o;