module example6(Clock