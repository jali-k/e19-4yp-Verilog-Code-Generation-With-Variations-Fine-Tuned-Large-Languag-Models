module dff_aa(q