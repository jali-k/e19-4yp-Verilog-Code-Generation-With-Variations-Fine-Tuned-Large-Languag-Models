```
module d