```SystemVerilog
// Create a module with one input and one output that behaves like a wire
module wire_assign(input in, output out);
    //assign out to in
    assign out = in;
endmodule
endmodule
```
### Result:
After running the test case, SystemVerilog Verific generates the following error:
```
>./vrun -v +acc +acc -p

vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:8: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:15: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:16: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:17: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:18: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:20: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:21: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:22: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:23: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:24: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:27: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:28: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:30: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:34: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:37: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:40: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:41: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:42: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:43: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:46: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:47: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:50: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:53: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:54: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:57: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:60: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:61: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:62: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:63: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:64: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:67: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:68: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:71: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:72: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:75: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:78: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:79: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:80: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:81: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:84: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:87: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:90: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:91: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:92: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:93: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:94: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:99: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:102: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:103: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:104: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:105: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:106: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:107: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:108: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:114: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:117: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:118: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:119: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:120: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:121: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:122: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:123: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:124: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:127: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:128: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14:131: vsim_verif: Error:.././/sv_lib/tb/tb_wire.sv:14: