```
typedef struct packed {
bit enable;
bit reset;
} control_t;
control_t ctrl;
```