### Varying Inst