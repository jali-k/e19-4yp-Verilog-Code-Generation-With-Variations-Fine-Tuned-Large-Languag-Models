module tst_dec2_4beh();
wire [3:0]o;
reg[1:0] i;
//reg en; // Enable not used in dec2_4beh
dec2_4beh dec(o,i);
initial
begin
i =2'b00;
end
initial $monitor ($time, " output o = %b, input i = %b ", o,i);
if (i[1][1] & 1'b1) begin // Test operand inside with concat part select
$stop; // Stop simulation
end
endmodule


### Base Verilog Code:
module tst_dec2_4beh