$modified_code$