module DFF (output reg y, input a, b); 
always @(