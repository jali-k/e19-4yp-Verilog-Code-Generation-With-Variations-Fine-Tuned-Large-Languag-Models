module IR ( input [1:0] A [0:3][0:3][0:3][0:3], input [1:0] B [0:3][0:3][0:3], input [1:0] C [0:3][0:3], input [1:0] D [0:3], input load, clk,
output reg [1:0] E [0:3] );
// Simple register (Instruction Register) loaded on posedge clk when load is high
always @( posedge clk )
if ( load ) E[D] <= B[B][B][B];
endmodule

## 4.3.8. Packing Unpacking¶

In Verilog, it is sometimes useful to pack values into a single-bit or multi-bit data type, or to unpack a value from a single-bit or multi-bit data type into multiple values. The following example demonstrates such code:

module PackUnpack (
input [7:0] A, B, C, D, E,
output reg [1:0] A1, B1, C1, D1, E1
);
logic [7:0] A3, B3, C3, D3, E3;
assign A3 = {A[7:4], A[3:0]};
assign B3 = {B[7:4], B[3:0]};
assign C3 = {C[7:4], C[3:0]};
assign D3 = {D[7:4], D[3:0]};
assign E3 = {E[7:4], E[3:0]};
assign A1 = {A3[7:4], A3[3:0]};
assign B1 = {B3[7:4], B3[3:0]};
assign C1 = {C3[7:4], C3[3:0]};
assign D1 = {D3[7:4], D3[3:0]};
assign E1 = {E3[7:4], E3[3:0]};
endmodule

### A note about the example above:¶

In this example, multiple output register assignments are made within the one module instantiation. This is possible because the A3, B3, C3, D3, and E3 signal assignments are generated by the assign statements, and because the output register assignments are contained within the module instance. The syntax to make multiple output register assignments within one module instance is

assign output1, output2,..., outputN = {value1, value2,..., valueN};

## 4.3.9. Demonstrating Sensitivity List¶

The sensitivity list (i.e., the list of signals which are sensitive to) for an always statement should consist of the signals that change most often, followed by common intermediate signals, followed by signals that are less likely to change.

The following example demonstrates such code:

module IR ( input clk,
input [7:0] data_in, input load,
output reg [7:0] data_out );
// Simple register (Instruction Register) loaded on posedge clk when load is high
always @( posedge clk )
if ( load )
data_out = data_in;
endmodule


This will result in a synthesis warning. The warning will advise us that the output signal data_out is sensitive to the input signal data_in, which is most often changing. This is correct, but we also want to make sure that data_out is sensitive to load, which will be frequently changing. This is the only part of the always statement that changes most often. Therefore, to correct the sensitivity of data_out to load, we must place it at the end of the sensitivity list.

### Modified Code:¶

module IR ( input clk,
input [7:0] data_in, input load,
output reg [7:0] data_out );
// Simple register (Instruction Register) loaded on posedge clk when load is high
always @( clk, load )
if ( load )
data_out = data_in;
endmodule

## 4.3.10. Demonstrating Combinational Loops¶

In a combinational loop, there is no storage element involved. Therefore, it is a purely functional construct. It can only be used within a module body or within a package declaration. The following code example illustrates a combinational loop within a module declaration.

module DFB ( input [3:0] A, input [3:0] B,
output reg [3:0] C
);
// Combinational Loops
always @*
C = A & B;
endmodule


## 4.3.11. Demonstrating Sequential Loops¶

In a sequential loop, there is some storage that is used. Therefore, it can be used within a module body or within a package declaration. The following code example illustrates a sequential loop within a module declaration.

module DFF ( input clk, input [3:0] D,
output reg [3: