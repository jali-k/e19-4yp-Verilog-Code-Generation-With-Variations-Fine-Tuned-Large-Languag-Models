module SchedDelayA (schedDelayA_inst);
wire clk;
wire rst;

reg [7:0] a, b;

schedDelayA_inst = @(posedge clk) begin
if (rst) a <= 1'b0;
a <= a + 1;
b <= a;
end
endmodule

How do you think it will change the generated verilog code? What is the impact on the circuit?

I am looking for answers that describe how this will change the generated verilog code in this particular case.

I have no idea how your compiler will treat it. It's not very likely to matter because it wouldn't add or change any functionality, but it's still wrong.

• The code I provided was generated by Lime. –  Apr 23 '20 at 22:16
• I am not sure what you are describing, but your schematic is correct. The first register input is just a wire. The second register input does not have a class handle, so it needs to be added and removed the same as a register. The second wire must also be created to be connected to the first register. –  Apr 23 '20 at 22:24
• Also, in your code, the third input is the reset. The class handle is used to define the third input in the verilog module. –  Apr 23 '20 at 22:27
• I am trying to understand what is the difference between the 1st and 3rd registers. What about the 2nd register? Are they the same? –  Apr 23 '20 at 22:31
• I used to think that the 1st and 3rd were the same, but I think they are separate registers. –  Apr 23 '20 at 22:36

The problem is that the code you have posted adds a third register, which has no class handle, to the module SchedDelayA. While the code will compile, and the resulting circuit will behave correctly, the code is incorrect. If you run the code through lint, the compiler will complain.

The code you have posted in the question is synthesized as follows, where:

• the first wire is a wire,
• the second wire is a reg[7:0]
• the third wire is a wire,

This is not a problem if the compiler creates the additional 3rd wire, but the code in the question is not synthesizable.

My understanding is that this is a bug in Lime, but I have no idea how it would handle this.

• The generated code for the schematic shows that the second wire is not a reg[7:0] but a wire. –  Apr 23 '20 at 22:19